module not_9b(in, out);

	input[8:0] in;
	output[8:0] out;

	assign out = ~(in);
endmodule
