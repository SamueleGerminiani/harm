module or_(out, a, b, c);

	input a,b,c;
	output out;

	assign out = a | b | c;
endmodule
