`timescale 1ns/1ps
module sin_lut(a, out);
	input  [31:0] a;
	output reg [31:0] out;
	wire   [10:0] index;

	always @(index)
	begin
		case(index)
			11'd0: out = 32'b00000000000000000000000001000000; // input=0.001953125, output=0.00195312375824
			11'd1: out = 32'b00000000000000000000000011000000; // input=0.005859375, output=0.00585934147244
			11'd2: out = 32'b00000000000000000000000101000000; // input=0.009765625, output=0.00976546978031
			11'd3: out = 32'b00000000000000000000000111000000; // input=0.013671875, output=0.0136714490791
			11'd4: out = 32'b00000000000000000000001001000000; // input=0.017578125, output=0.0175772197684
			11'd5: out = 32'b00000000000000000000001011000000; // input=0.021484375, output=0.021482722251
			11'd6: out = 32'b00000000000000000000001101000000; // input=0.025390625, output=0.0253878969337
			11'd7: out = 32'b00000000000000000000001111000000; // input=0.029296875, output=0.0292926842283
			11'd8: out = 32'b00000000000000000000010001000000; // input=0.033203125, output=0.0331970245525
			11'd9: out = 32'b00000000000000000000010011000000; // input=0.037109375, output=0.0371008583311
			11'd10: out = 32'b00000000000000000000010101000000; // input=0.041015625, output=0.0410041259961
			11'd11: out = 32'b00000000000000000000010111000000; // input=0.044921875, output=0.0449067679887
			11'd12: out = 32'b00000000000000000000011000111111; // input=0.048828125, output=0.0488087247592
			11'd13: out = 32'b00000000000000000000011010111111; // input=0.052734375, output=0.0527099367686
			11'd14: out = 32'b00000000000000000000011100111111; // input=0.056640625, output=0.0566103444893
			11'd15: out = 32'b00000000000000000000011110111111; // input=0.060546875, output=0.0605098884057
			11'd16: out = 32'b00000000000000000000100000111111; // input=0.064453125, output=0.0644085090157
			11'd17: out = 32'b00000000000000000000100010111110; // input=0.068359375, output=0.0683061468311
			11'd18: out = 32'b00000000000000000000100100111110; // input=0.072265625, output=0.0722027423787
			11'd19: out = 32'b00000000000000000000100110111110; // input=0.076171875, output=0.0760982362014
			11'd20: out = 32'b00000000000000000000101000111101; // input=0.080078125, output=0.0799925688585
			11'd21: out = 32'b00000000000000000000101010111101; // input=0.083984375, output=0.0838856809275
			11'd22: out = 32'b00000000000000000000101100111100; // input=0.087890625, output=0.0877775130042
			11'd23: out = 32'b00000000000000000000101110111100; // input=0.091796875, output=0.091668005704
			11'd24: out = 32'b00000000000000000000110000111011; // input=0.095703125, output=0.0955570996629
			11'd25: out = 32'b00000000000000000000110010111011; // input=0.099609375, output=0.099444735538
			11'd26: out = 32'b00000000000000000000110100111010; // input=0.103515625, output=0.103330854009
			11'd27: out = 32'b00000000000000000000110110111001; // input=0.107421875, output=0.107215395778
			11'd28: out = 32'b00000000000000000000111000111000; // input=0.111328125, output=0.111098301572
			11'd29: out = 32'b00000000000000000000111010111000; // input=0.115234375, output=0.114979512142
			11'd30: out = 32'b00000000000000000000111100110111; // input=0.119140625, output=0.118858968267
			11'd31: out = 32'b00000000000000000000111110110110; // input=0.123046875, output=0.12273661075
			11'd32: out = 32'b00000000000000000001000000110101; // input=0.126953125, output=0.126612380424
			11'd33: out = 32'b00000000000000000001000010110100; // input=0.130859375, output=0.130486218148
			11'd34: out = 32'b00000000000000000001000100110011; // input=0.134765625, output=0.134358064813
			11'd35: out = 32'b00000000000000000001000110110001; // input=0.138671875, output=0.13822786134
			11'd36: out = 32'b00000000000000000001001000110000; // input=0.142578125, output=0.142095548679
			11'd37: out = 32'b00000000000000000001001010101111; // input=0.146484375, output=0.145961067815
			11'd38: out = 32'b00000000000000000001001100101101; // input=0.150390625, output=0.149824359765
			11'd39: out = 32'b00000000000000000001001110101100; // input=0.154296875, output=0.153685365579
			11'd40: out = 32'b00000000000000000001010000101010; // input=0.158203125, output=0.157544026344
			11'd41: out = 32'b00000000000000000001010010101001; // input=0.162109375, output=0.161400283181
			11'd42: out = 32'b00000000000000000001010100100111; // input=0.166015625, output=0.165254077248
			11'd43: out = 32'b00000000000000000001010110100101; // input=0.169921875, output=0.169105349741
			11'd44: out = 32'b00000000000000000001011000100011; // input=0.173828125, output=0.172954041894
			11'd45: out = 32'b00000000000000000001011010100001; // input=0.177734375, output=0.176800094982
			11'd46: out = 32'b00000000000000000001011100011111; // input=0.181640625, output=0.180643450318
			11'd47: out = 32'b00000000000000000001011110011101; // input=0.185546875, output=0.184484049257
			11'd48: out = 32'b00000000000000000001100000011011; // input=0.189453125, output=0.188321833196
			11'd49: out = 32'b00000000000000000001100010011001; // input=0.193359375, output=0.192156743576
			11'd50: out = 32'b00000000000000000001100100010110; // input=0.197265625, output=0.19598872188
			11'd51: out = 32'b00000000000000000001100110010100; // input=0.201171875, output=0.199817709638
			11'd52: out = 32'b00000000000000000001101000010001; // input=0.205078125, output=0.203643648423
			11'd53: out = 32'b00000000000000000001101010001110; // input=0.208984375, output=0.207466479857
			11'd54: out = 32'b00000000000000000001101100001011; // input=0.212890625, output=0.211286145607
			11'd55: out = 32'b00000000000000000001101110001000; // input=0.216796875, output=0.215102587391
			11'd56: out = 32'b00000000000000000001110000000101; // input=0.220703125, output=0.218915746974
			11'd57: out = 32'b00000000000000000001110010000010; // input=0.224609375, output=0.222725566172
			11'd58: out = 32'b00000000000000000001110011111111; // input=0.228515625, output=0.226531986852
			11'd59: out = 32'b00000000000000000001110101111100; // input=0.232421875, output=0.230334950932
			11'd60: out = 32'b00000000000000000001110111111000; // input=0.236328125, output=0.234134400385
			11'd61: out = 32'b00000000000000000001111001110100; // input=0.240234375, output=0.237930277234
			11'd62: out = 32'b00000000000000000001111011110001; // input=0.244140625, output=0.241722523561
			11'd63: out = 32'b00000000000000000001111101101101; // input=0.248046875, output=0.245511081499
			11'd64: out = 32'b00000000000000000001111111101001; // input=0.251953125, output=0.24929589324
			11'd65: out = 32'b00000000000000000010000001100101; // input=0.255859375, output=0.253076901032
			11'd66: out = 32'b00000000000000000010000011100001; // input=0.259765625, output=0.256854047182
			11'd67: out = 32'b00000000000000000010000101011100; // input=0.263671875, output=0.260627274056
			11'd68: out = 32'b00000000000000000010000111011000; // input=0.267578125, output=0.264396524078
			11'd69: out = 32'b00000000000000000010001001010011; // input=0.271484375, output=0.268161739734
			11'd70: out = 32'b00000000000000000010001011001110; // input=0.275390625, output=0.271922863572
			11'd71: out = 32'b00000000000000000010001101001001; // input=0.279296875, output=0.275679838202
			11'd72: out = 32'b00000000000000000010001111000100; // input=0.283203125, output=0.279432606296
			11'd73: out = 32'b00000000000000000010010000111111; // input=0.287109375, output=0.283181110593
			11'd74: out = 32'b00000000000000000010010010111010; // input=0.291015625, output=0.286925293895
			11'd75: out = 32'b00000000000000000010010100110101; // input=0.294921875, output=0.290665099069
			11'd76: out = 32'b00000000000000000010010110101111; // input=0.298828125, output=0.294400469052
			11'd77: out = 32'b00000000000000000010011000101001; // input=0.302734375, output=0.298131346846
			11'd78: out = 32'b00000000000000000010011010100011; // input=0.306640625, output=0.301857675522
			11'd79: out = 32'b00000000000000000010011100011101; // input=0.310546875, output=0.305579398221
			11'd80: out = 32'b00000000000000000010011110010111; // input=0.314453125, output=0.309296458155
			11'd81: out = 32'b00000000000000000010100000010001; // input=0.318359375, output=0.313008798605
			11'd82: out = 32'b00000000000000000010100010001010; // input=0.322265625, output=0.316716362927
			11'd83: out = 32'b00000000000000000010100100000011; // input=0.326171875, output=0.320419094546
			11'd84: out = 32'b00000000000000000010100101111101; // input=0.330078125, output=0.324116936964
			11'd85: out = 32'b00000000000000000010100111110110; // input=0.333984375, output=0.327809833756
			11'd86: out = 32'b00000000000000000010101001101111; // input=0.337890625, output=0.331497728574
			11'd87: out = 32'b00000000000000000010101011100111; // input=0.341796875, output=0.335180565144
			11'd88: out = 32'b00000000000000000010101101100000; // input=0.345703125, output=0.338858287271
			11'd89: out = 32'b00000000000000000010101111011000; // input=0.349609375, output=0.342530838838
			11'd90: out = 32'b00000000000000000010110001010000; // input=0.353515625, output=0.346198163805
			11'd91: out = 32'b00000000000000000010110011001000; // input=0.357421875, output=0.349860206215
			11'd92: out = 32'b00000000000000000010110101000000; // input=0.361328125, output=0.353516910188
			11'd93: out = 32'b00000000000000000010110110111000; // input=0.365234375, output=0.357168219928
			11'd94: out = 32'b00000000000000000010111000101111; // input=0.369140625, output=0.36081407972
			11'd95: out = 32'b00000000000000000010111010100110; // input=0.373046875, output=0.364454433933
			11'd96: out = 32'b00000000000000000010111100011110; // input=0.376953125, output=0.36808922702
			11'd97: out = 32'b00000000000000000010111110010100; // input=0.380859375, output=0.371718403519
			11'd98: out = 32'b00000000000000000011000000001011; // input=0.384765625, output=0.375341908052
			11'd99: out = 32'b00000000000000000011000010000010; // input=0.388671875, output=0.378959685329
			11'd100: out = 32'b00000000000000000011000011111000; // input=0.392578125, output=0.382571680148
			11'd101: out = 32'b00000000000000000011000101101110; // input=0.396484375, output=0.386177837393
			11'd102: out = 32'b00000000000000000011000111100100; // input=0.400390625, output=0.38977810204
			11'd103: out = 32'b00000000000000000011001001011010; // input=0.404296875, output=0.393372419153
			11'd104: out = 32'b00000000000000000011001011010000; // input=0.408203125, output=0.396960733886
			11'd105: out = 32'b00000000000000000011001101000101; // input=0.412109375, output=0.400542991487
			11'd106: out = 32'b00000000000000000011001110111010; // input=0.416015625, output=0.404119137295
			11'd107: out = 32'b00000000000000000011010000101111; // input=0.419921875, output=0.407689116742
			11'd108: out = 32'b00000000000000000011010010100100; // input=0.423828125, output=0.411252875354
			11'd109: out = 32'b00000000000000000011010100011001; // input=0.427734375, output=0.414810358754
			11'd110: out = 32'b00000000000000000011010110001101; // input=0.431640625, output=0.418361512658
			11'd111: out = 32'b00000000000000000011011000000001; // input=0.435546875, output=0.42190628288
			11'd112: out = 32'b00000000000000000011011001110101; // input=0.439453125, output=0.425444615332
			11'd113: out = 32'b00000000000000000011011011101001; // input=0.443359375, output=0.428976456021
			11'd114: out = 32'b00000000000000000011011101011100; // input=0.447265625, output=0.432501751058
			11'd115: out = 32'b00000000000000000011011111010000; // input=0.451171875, output=0.436020446651
			11'd116: out = 32'b00000000000000000011100001000011; // input=0.455078125, output=0.439532489107
			11'd117: out = 32'b00000000000000000011100010110101; // input=0.458984375, output=0.443037824839
			11'd118: out = 32'b00000000000000000011100100101000; // input=0.462890625, output=0.446536400359
			11'd119: out = 32'b00000000000000000011100110011011; // input=0.466796875, output=0.450028162283
			11'd120: out = 32'b00000000000000000011101000001101; // input=0.470703125, output=0.45351305733
			11'd121: out = 32'b00000000000000000011101001111111; // input=0.474609375, output=0.456991032326
			11'd122: out = 32'b00000000000000000011101011110000; // input=0.478515625, output=0.460462034202
			11'd123: out = 32'b00000000000000000011101101100010; // input=0.482421875, output=0.463926009993
			11'd124: out = 32'b00000000000000000011101111010011; // input=0.486328125, output=0.467382906844
			11'd125: out = 32'b00000000000000000011110001000100; // input=0.490234375, output=0.470832672007
			11'd126: out = 32'b00000000000000000011110010110101; // input=0.494140625, output=0.474275252843
			11'd127: out = 32'b00000000000000000011110100100110; // input=0.498046875, output=0.477710596821
			11'd128: out = 32'b00000000000000000011110110010110; // input=0.501953125, output=0.481138651524
			11'd129: out = 32'b00000000000000000011111000000110; // input=0.505859375, output=0.484559364643
			11'd130: out = 32'b00000000000000000011111001110110; // input=0.509765625, output=0.487972683983
			11'd131: out = 32'b00000000000000000011111011100101; // input=0.513671875, output=0.491378557459
			11'd132: out = 32'b00000000000000000011111101010101; // input=0.517578125, output=0.494776933103
			11'd133: out = 32'b00000000000000000011111111000100; // input=0.521484375, output=0.49816775906
			11'd134: out = 32'b00000000000000000100000000110011; // input=0.525390625, output=0.50155098359
			11'd135: out = 32'b00000000000000000100000010100001; // input=0.529296875, output=0.504926555069
			11'd136: out = 32'b00000000000000000100000100010000; // input=0.533203125, output=0.50829442199
			11'd137: out = 32'b00000000000000000100000101111110; // input=0.537109375, output=0.511654532964
			11'd138: out = 32'b00000000000000000100000111101100; // input=0.541015625, output=0.515006836719
			11'd139: out = 32'b00000000000000000100001001011001; // input=0.544921875, output=0.518351282103
			11'd140: out = 32'b00000000000000000100001011000111; // input=0.548828125, output=0.521687818084
			11'd141: out = 32'b00000000000000000100001100110100; // input=0.552734375, output=0.525016393751
			11'd142: out = 32'b00000000000000000100001110100001; // input=0.556640625, output=0.528336958314
			11'd143: out = 32'b00000000000000000100010000001101; // input=0.560546875, output=0.531649461105
			11'd144: out = 32'b00000000000000000100010001111001; // input=0.564453125, output=0.534953851579
			11'd145: out = 32'b00000000000000000100010011100101; // input=0.568359375, output=0.538250079316
			11'd146: out = 32'b00000000000000000100010101010001; // input=0.572265625, output=0.541538094019
			11'd147: out = 32'b00000000000000000100010110111101; // input=0.576171875, output=0.544817845516
			11'd148: out = 32'b00000000000000000100011000101000; // input=0.580078125, output=0.548089283764
			11'd149: out = 32'b00000000000000000100011010010011; // input=0.583984375, output=0.551352358843
			11'd150: out = 32'b00000000000000000100011011111101; // input=0.587890625, output=0.554607020964
			11'd151: out = 32'b00000000000000000100011101101000; // input=0.591796875, output=0.557853220464
			11'd152: out = 32'b00000000000000000100011111010010; // input=0.595703125, output=0.561090907811
			11'd153: out = 32'b00000000000000000100100000111100; // input=0.599609375, output=0.5643200336
			11'd154: out = 32'b00000000000000000100100010100101; // input=0.603515625, output=0.56754054856
			11'd155: out = 32'b00000000000000000100100100001110; // input=0.607421875, output=0.570752403549
			11'd156: out = 32'b00000000000000000100100101110111; // input=0.611328125, output=0.573955549559
			11'd157: out = 32'b00000000000000000100100111100000; // input=0.615234375, output=0.577149937714
			11'd158: out = 32'b00000000000000000100101001001000; // input=0.619140625, output=0.58033551927
			11'd159: out = 32'b00000000000000000100101010110001; // input=0.623046875, output=0.583512245621
			11'd160: out = 32'b00000000000000000100101100011000; // input=0.626953125, output=0.586680068292
			11'd161: out = 32'b00000000000000000100101110000000; // input=0.630859375, output=0.589838938948
			11'd162: out = 32'b00000000000000000100101111100111; // input=0.634765625, output=0.592988809387
			11'd163: out = 32'b00000000000000000100110001001110; // input=0.638671875, output=0.596129631546
			11'd164: out = 32'b00000000000000000100110010110101; // input=0.642578125, output=0.599261357501
			11'd165: out = 32'b00000000000000000100110100011011; // input=0.646484375, output=0.602383939464
			11'd166: out = 32'b00000000000000000100110110000001; // input=0.650390625, output=0.60549732979
			11'd167: out = 32'b00000000000000000100110111100111; // input=0.654296875, output=0.608601480971
			11'd168: out = 32'b00000000000000000100111001001100; // input=0.658203125, output=0.611696345643
			11'd169: out = 32'b00000000000000000100111010110001; // input=0.662109375, output=0.614781876581
			11'd170: out = 32'b00000000000000000100111100010110; // input=0.666015625, output=0.617858026704
			11'd171: out = 32'b00000000000000000100111101111010; // input=0.669921875, output=0.620924749074
			11'd172: out = 32'b00000000000000000100111111011111; // input=0.673828125, output=0.623981996896
			11'd173: out = 32'b00000000000000000101000001000011; // input=0.677734375, output=0.62702972352
			11'd174: out = 32'b00000000000000000101000010100110; // input=0.681640625, output=0.630067882443
			11'd175: out = 32'b00000000000000000101000100001001; // input=0.685546875, output=0.633096427304
			11'd176: out = 32'b00000000000000000101000101101100; // input=0.689453125, output=0.636115311893
			11'd177: out = 32'b00000000000000000101000111001111; // input=0.693359375, output=0.639124490145
			11'd178: out = 32'b00000000000000000101001000110001; // input=0.697265625, output=0.642123916144
			11'd179: out = 32'b00000000000000000101001010010011; // input=0.701171875, output=0.645113544122
			11'd180: out = 32'b00000000000000000101001011110101; // input=0.705078125, output=0.64809332846
			11'd181: out = 32'b00000000000000000101001101010110; // input=0.708984375, output=0.651063223692
			11'd182: out = 32'b00000000000000000101001110110111; // input=0.712890625, output=0.6540231845
			11'd183: out = 32'b00000000000000000101010000011000; // input=0.716796875, output=0.65697316572
			11'd184: out = 32'b00000000000000000101010001111000; // input=0.720703125, output=0.659913122336
			11'd185: out = 32'b00000000000000000101010011011000; // input=0.724609375, output=0.662843009491
			11'd186: out = 32'b00000000000000000101010100111000; // input=0.728515625, output=0.665762782477
			11'd187: out = 32'b00000000000000000101010110010111; // input=0.732421875, output=0.668672396741
			11'd188: out = 32'b00000000000000000101010111110110; // input=0.736328125, output=0.671571807888
			11'd189: out = 32'b00000000000000000101011001010101; // input=0.740234375, output=0.674460971675
			11'd190: out = 32'b00000000000000000101011010110011; // input=0.744140625, output=0.677339844018
			11'd191: out = 32'b00000000000000000101011100010001; // input=0.748046875, output=0.680208380988
			11'd192: out = 32'b00000000000000000101011101101111; // input=0.751953125, output=0.683066538814
			11'd193: out = 32'b00000000000000000101011111001100; // input=0.755859375, output=0.685914273886
			11'd194: out = 32'b00000000000000000101100000101001; // input=0.759765625, output=0.68875154275
			11'd195: out = 32'b00000000000000000101100010000110; // input=0.763671875, output=0.691578302113
			11'd196: out = 32'b00000000000000000101100011100010; // input=0.767578125, output=0.694394508842
			11'd197: out = 32'b00000000000000000101100100111110; // input=0.771484375, output=0.697200119965
			11'd198: out = 32'b00000000000000000101100110011001; // input=0.775390625, output=0.699995092672
			11'd199: out = 32'b00000000000000000101100111110101; // input=0.779296875, output=0.702779384315
			11'd200: out = 32'b00000000000000000101101001010000; // input=0.783203125, output=0.705552952409
			11'd201: out = 32'b00000000000000000101101010101010; // input=0.787109375, output=0.708315754633
			11'd202: out = 32'b00000000000000000101101100000100; // input=0.791015625, output=0.711067748831
			11'd203: out = 32'b00000000000000000101101101011110; // input=0.794921875, output=0.713808893009
			11'd204: out = 32'b00000000000000000101101110111000; // input=0.798828125, output=0.716539145342
			11'd205: out = 32'b00000000000000000101110000010001; // input=0.802734375, output=0.719258464169
			11'd206: out = 32'b00000000000000000101110001101001; // input=0.806640625, output=0.721966807997
			11'd207: out = 32'b00000000000000000101110011000010; // input=0.810546875, output=0.7246641355
			11'd208: out = 32'b00000000000000000101110100011010; // input=0.814453125, output=0.727350405519
			11'd209: out = 32'b00000000000000000101110101110001; // input=0.818359375, output=0.730025577067
			11'd210: out = 32'b00000000000000000101110111001001; // input=0.822265625, output=0.732689609322
			11'd211: out = 32'b00000000000000000101111000100000; // input=0.826171875, output=0.735342461635
			11'd212: out = 32'b00000000000000000101111001110110; // input=0.830078125, output=0.737984093527
			11'd213: out = 32'b00000000000000000101111011001100; // input=0.833984375, output=0.740614464689
			11'd214: out = 32'b00000000000000000101111100100010; // input=0.837890625, output=0.743233534986
			11'd215: out = 32'b00000000000000000101111101111000; // input=0.841796875, output=0.745841264454
			11'd216: out = 32'b00000000000000000101111111001101; // input=0.845703125, output=0.748437613302
			11'd217: out = 32'b00000000000000000110000000100010; // input=0.849609375, output=0.751022541912
			11'd218: out = 32'b00000000000000000110000001110110; // input=0.853515625, output=0.753596010843
			11'd219: out = 32'b00000000000000000110000011001010; // input=0.857421875, output=0.756157980826
			11'd220: out = 32'b00000000000000000110000100011101; // input=0.861328125, output=0.758708412768
			11'd221: out = 32'b00000000000000000110000101110001; // input=0.865234375, output=0.761247267753
			11'd222: out = 32'b00000000000000000110000111000011; // input=0.869140625, output=0.763774507042
			11'd223: out = 32'b00000000000000000110001000010110; // input=0.873046875, output=0.766290092071
			11'd224: out = 32'b00000000000000000110001001101000; // input=0.876953125, output=0.768793984456
			11'd225: out = 32'b00000000000000000110001010111010; // input=0.880859375, output=0.771286145991
			11'd226: out = 32'b00000000000000000110001100001011; // input=0.884765625, output=0.773766538648
			11'd227: out = 32'b00000000000000000110001101011100; // input=0.888671875, output=0.77623512458
			11'd228: out = 32'b00000000000000000110001110101100; // input=0.892578125, output=0.778691866119
			11'd229: out = 32'b00000000000000000110001111111100; // input=0.896484375, output=0.781136725778
			11'd230: out = 32'b00000000000000000110010001001100; // input=0.900390625, output=0.783569666252
			11'd231: out = 32'b00000000000000000110010010011011; // input=0.904296875, output=0.785990650417
			11'd232: out = 32'b00000000000000000110010011101010; // input=0.908203125, output=0.788399641331
			11'd233: out = 32'b00000000000000000110010100111001; // input=0.912109375, output=0.790796602237
			11'd234: out = 32'b00000000000000000110010110000111; // input=0.916015625, output=0.79318149656
			11'd235: out = 32'b00000000000000000110010111010101; // input=0.919921875, output=0.795554287909
			11'd236: out = 32'b00000000000000000110011000100010; // input=0.923828125, output=0.797914940078
			11'd237: out = 32'b00000000000000000110011001101111; // input=0.927734375, output=0.800263417047
			11'd238: out = 32'b00000000000000000110011010111100; // input=0.931640625, output=0.802599682981
			11'd239: out = 32'b00000000000000000110011100001000; // input=0.935546875, output=0.804923702231
			11'd240: out = 32'b00000000000000000110011101010011; // input=0.939453125, output=0.807235439336
			11'd241: out = 32'b00000000000000000110011110011111; // input=0.943359375, output=0.809534859021
			11'd242: out = 32'b00000000000000000110011111101010; // input=0.947265625, output=0.8118219262
			11'd243: out = 32'b00000000000000000110100000110100; // input=0.951171875, output=0.814096605976
			11'd244: out = 32'b00000000000000000110100001111110; // input=0.955078125, output=0.816358863639
			11'd245: out = 32'b00000000000000000110100011001000; // input=0.958984375, output=0.81860866467
			11'd246: out = 32'b00000000000000000110100100010001; // input=0.962890625, output=0.82084597474
			11'd247: out = 32'b00000000000000000110100101011010; // input=0.966796875, output=0.82307075971
			11'd248: out = 32'b00000000000000000110100110100011; // input=0.970703125, output=0.825282985633
			11'd249: out = 32'b00000000000000000110100111101011; // input=0.974609375, output=0.827482618753
			11'd250: out = 32'b00000000000000000110101000110011; // input=0.978515625, output=0.829669625507
			11'd251: out = 32'b00000000000000000110101001111010; // input=0.982421875, output=0.831843972523
			11'd252: out = 32'b00000000000000000110101011000001; // input=0.986328125, output=0.834005626623
			11'd253: out = 32'b00000000000000000110101100000111; // input=0.990234375, output=0.836154554823
			11'd254: out = 32'b00000000000000000110101101001101; // input=0.994140625, output=0.838290724334
			11'd255: out = 32'b00000000000000000110101110010011; // input=0.998046875, output=0.84041410256
			11'd256: out = 32'b00000000000000000110101111011000; // input=1.001953125, output=0.8425246571
			11'd257: out = 32'b00000000000000000110110000011101; // input=1.005859375, output=0.844622355751
			11'd258: out = 32'b00000000000000000110110001100001; // input=1.009765625, output=0.846707166504
			11'd259: out = 32'b00000000000000000110110010100101; // input=1.013671875, output=0.848779057547
			11'd260: out = 32'b00000000000000000110110011101000; // input=1.017578125, output=0.850837997266
			11'd261: out = 32'b00000000000000000110110100101011; // input=1.021484375, output=0.852883954244
			11'd262: out = 32'b00000000000000000110110101101110; // input=1.025390625, output=0.854916897262
			11'd263: out = 32'b00000000000000000110110110110000; // input=1.029296875, output=0.8569367953
			11'd264: out = 32'b00000000000000000110110111110010; // input=1.033203125, output=0.858943617537
			11'd265: out = 32'b00000000000000000110111000110011; // input=1.037109375, output=0.860937333352
			11'd266: out = 32'b00000000000000000110111001110100; // input=1.041015625, output=0.862917912321
			11'd267: out = 32'b00000000000000000110111010110101; // input=1.044921875, output=0.864885324225
			11'd268: out = 32'b00000000000000000110111011110101; // input=1.048828125, output=0.866839539044
			11'd269: out = 32'b00000000000000000110111100110100; // input=1.052734375, output=0.868780526957
			11'd270: out = 32'b00000000000000000110111101110011; // input=1.056640625, output=0.870708258348
			11'd271: out = 32'b00000000000000000110111110110010; // input=1.060546875, output=0.872622703803
			11'd272: out = 32'b00000000000000000110111111110000; // input=1.064453125, output=0.874523834109
			11'd273: out = 32'b00000000000000000111000000101110; // input=1.068359375, output=0.876411620257
			11'd274: out = 32'b00000000000000000111000001101100; // input=1.072265625, output=0.878286033441
			11'd275: out = 32'b00000000000000000111000010101001; // input=1.076171875, output=0.880147045062
			11'd276: out = 32'b00000000000000000111000011100101; // input=1.080078125, output=0.881994626722
			11'd277: out = 32'b00000000000000000111000100100001; // input=1.083984375, output=0.883828750229
			11'd278: out = 32'b00000000000000000111000101011101; // input=1.087890625, output=0.885649387596
			11'd279: out = 32'b00000000000000000111000110011000; // input=1.091796875, output=0.887456511044
			11'd280: out = 32'b00000000000000000111000111010011; // input=1.095703125, output=0.889250092997
			11'd281: out = 32'b00000000000000000111001000001101; // input=1.099609375, output=0.891030106087
			11'd282: out = 32'b00000000000000000111001001000111; // input=1.103515625, output=0.892796523155
			11'd283: out = 32'b00000000000000000111001010000001; // input=1.107421875, output=0.894549317246
			11'd284: out = 32'b00000000000000000111001010111010; // input=1.111328125, output=0.896288461615
			11'd285: out = 32'b00000000000000000111001011110010; // input=1.115234375, output=0.898013929725
			11'd286: out = 32'b00000000000000000111001100101010; // input=1.119140625, output=0.899725695247
			11'd287: out = 32'b00000000000000000111001101100010; // input=1.123046875, output=0.901423732062
			11'd288: out = 32'b00000000000000000111001110011001; // input=1.126953125, output=0.90310801426
			11'd289: out = 32'b00000000000000000111001111010000; // input=1.130859375, output=0.90477851614
			11'd290: out = 32'b00000000000000000111010000000110; // input=1.134765625, output=0.906435212214
			11'd291: out = 32'b00000000000000000111010000111100; // input=1.138671875, output=0.908078077202
			11'd292: out = 32'b00000000000000000111010001110001; // input=1.142578125, output=0.909707086035
			11'd293: out = 32'b00000000000000000111010010100110; // input=1.146484375, output=0.911322213858
			11'd294: out = 32'b00000000000000000111010011011011; // input=1.150390625, output=0.912923436025
			11'd295: out = 32'b00000000000000000111010100001111; // input=1.154296875, output=0.914510728103
			11'd296: out = 32'b00000000000000000111010101000010; // input=1.158203125, output=0.916084065873
			11'd297: out = 32'b00000000000000000111010101110101; // input=1.162109375, output=0.917643425327
			11'd298: out = 32'b00000000000000000111010110101000; // input=1.166015625, output=0.919188782671
			11'd299: out = 32'b00000000000000000111010111011010; // input=1.169921875, output=0.920720114326
			11'd300: out = 32'b00000000000000000111011000001100; // input=1.173828125, output=0.922237396924
			11'd301: out = 32'b00000000000000000111011000111101; // input=1.177734375, output=0.923740607315
			11'd302: out = 32'b00000000000000000111011001101110; // input=1.181640625, output=0.92522972256
			11'd303: out = 32'b00000000000000000111011010011110; // input=1.185546875, output=0.926704719938
			11'd304: out = 32'b00000000000000000111011011001110; // input=1.189453125, output=0.928165576942
			11'd305: out = 32'b00000000000000000111011011111110; // input=1.193359375, output=0.929612271281
			11'd306: out = 32'b00000000000000000111011100101100; // input=1.197265625, output=0.931044780881
			11'd307: out = 32'b00000000000000000111011101011011; // input=1.201171875, output=0.932463083883
			11'd308: out = 32'b00000000000000000111011110001001; // input=1.205078125, output=0.933867158646
			11'd309: out = 32'b00000000000000000111011110110111; // input=1.208984375, output=0.935256983744
			11'd310: out = 32'b00000000000000000111011111100100; // input=1.212890625, output=0.936632537972
			11'd311: out = 32'b00000000000000000111100000010000; // input=1.216796875, output=0.93799380034
			11'd312: out = 32'b00000000000000000111100000111100; // input=1.220703125, output=0.939340750076
			11'd313: out = 32'b00000000000000000111100001101000; // input=1.224609375, output=0.940673366629
			11'd314: out = 32'b00000000000000000111100010010011; // input=1.228515625, output=0.941991629663
			11'd315: out = 32'b00000000000000000111100010111110; // input=1.232421875, output=0.943295519063
			11'd316: out = 32'b00000000000000000111100011101000; // input=1.236328125, output=0.944585014935
			11'd317: out = 32'b00000000000000000111100100010010; // input=1.240234375, output=0.945860097601
			11'd318: out = 32'b00000000000000000111100100111011; // input=1.244140625, output=0.947120747606
			11'd319: out = 32'b00000000000000000111100101100100; // input=1.248046875, output=0.948366945714
			11'd320: out = 32'b00000000000000000111100110001100; // input=1.251953125, output=0.949598672909
			11'd321: out = 32'b00000000000000000111100110110100; // input=1.255859375, output=0.950815910397
			11'd322: out = 32'b00000000000000000111100111011100; // input=1.259765625, output=0.952018639603
			11'd323: out = 32'b00000000000000000111101000000011; // input=1.263671875, output=0.953206842177
			11'd324: out = 32'b00000000000000000111101000101001; // input=1.267578125, output=0.954380499987
			11'd325: out = 32'b00000000000000000111101001001111; // input=1.271484375, output=0.955539595124
			11'd326: out = 32'b00000000000000000111101001110101; // input=1.275390625, output=0.956684109903
			11'd327: out = 32'b00000000000000000111101010011010; // input=1.279296875, output=0.95781402686
			11'd328: out = 32'b00000000000000000111101010111110; // input=1.283203125, output=0.958929328753
			11'd329: out = 32'b00000000000000000111101011100010; // input=1.287109375, output=0.960029998564
			11'd330: out = 32'b00000000000000000111101100000110; // input=1.291015625, output=0.961116019499
			11'd331: out = 32'b00000000000000000111101100101001; // input=1.294921875, output=0.962187374985
			11'd332: out = 32'b00000000000000000111101101001100; // input=1.298828125, output=0.963244048676
			11'd333: out = 32'b00000000000000000111101101101110; // input=1.302734375, output=0.964286024448
			11'd334: out = 32'b00000000000000000111101110001111; // input=1.306640625, output=0.965313286402
			11'd335: out = 32'b00000000000000000111101110110001; // input=1.310546875, output=0.966325818863
			11'd336: out = 32'b00000000000000000111101111010001; // input=1.314453125, output=0.96732360638
			11'd337: out = 32'b00000000000000000111101111110001; // input=1.318359375, output=0.96830663373
			11'd338: out = 32'b00000000000000000111110000010001; // input=1.322265625, output=0.969274885911
			11'd339: out = 32'b00000000000000000111110000110000; // input=1.326171875, output=0.970228348151
			11'd340: out = 32'b00000000000000000111110001001111; // input=1.330078125, output=0.971167005899
			11'd341: out = 32'b00000000000000000111110001101101; // input=1.333984375, output=0.972090844834
			11'd342: out = 32'b00000000000000000111110010001011; // input=1.337890625, output=0.972999850858
			11'd343: out = 32'b00000000000000000111110010101001; // input=1.341796875, output=0.973894010102
			11'd344: out = 32'b00000000000000000111110011000101; // input=1.345703125, output=0.974773308922
			11'd345: out = 32'b00000000000000000111110011100010; // input=1.349609375, output=0.9756377339
			11'd346: out = 32'b00000000000000000111110011111110; // input=1.353515625, output=0.976487271847
			11'd347: out = 32'b00000000000000000111110100011001; // input=1.357421875, output=0.977321909799
			11'd348: out = 32'b00000000000000000111110100110100; // input=1.361328125, output=0.978141635021
			11'd349: out = 32'b00000000000000000111110101001110; // input=1.365234375, output=0.978946435006
			11'd350: out = 32'b00000000000000000111110101101000; // input=1.369140625, output=0.979736297472
			11'd351: out = 32'b00000000000000000111110110000001; // input=1.373046875, output=0.980511210368
			11'd352: out = 32'b00000000000000000111110110011010; // input=1.376953125, output=0.981271161869
			11'd353: out = 32'b00000000000000000111110110110011; // input=1.380859375, output=0.98201614038
			11'd354: out = 32'b00000000000000000111110111001011; // input=1.384765625, output=0.982746134532
			11'd355: out = 32'b00000000000000000111110111100010; // input=1.388671875, output=0.983461133188
			11'd356: out = 32'b00000000000000000111110111111001; // input=1.392578125, output=0.984161125436
			11'd357: out = 32'b00000000000000000111111000001111; // input=1.396484375, output=0.984846100597
			11'd358: out = 32'b00000000000000000111111000100101; // input=1.400390625, output=0.985516048218
			11'd359: out = 32'b00000000000000000111111000111011; // input=1.404296875, output=0.986170958077
			11'd360: out = 32'b00000000000000000111111001010000; // input=1.408203125, output=0.98681082018
			11'd361: out = 32'b00000000000000000111111001100100; // input=1.412109375, output=0.987435624764
			11'd362: out = 32'b00000000000000000111111001111000; // input=1.416015625, output=0.988045362295
			11'd363: out = 32'b00000000000000000111111010001100; // input=1.419921875, output=0.98864002347
			11'd364: out = 32'b00000000000000000111111010011111; // input=1.423828125, output=0.989219599214
			11'd365: out = 32'b00000000000000000111111010110001; // input=1.427734375, output=0.989784080684
			11'd366: out = 32'b00000000000000000111111011000011; // input=1.431640625, output=0.990333459267
			11'd367: out = 32'b00000000000000000111111011010101; // input=1.435546875, output=0.99086772658
			11'd368: out = 32'b00000000000000000111111011100110; // input=1.439453125, output=0.991386874471
			11'd369: out = 32'b00000000000000000111111011110110; // input=1.443359375, output=0.991890895017
			11'd370: out = 32'b00000000000000000111111100000110; // input=1.447265625, output=0.992379780529
			11'd371: out = 32'b00000000000000000111111100010110; // input=1.451171875, output=0.992853523546
			11'd372: out = 32'b00000000000000000111111100100101; // input=1.455078125, output=0.99331211684
			11'd373: out = 32'b00000000000000000111111100110011; // input=1.458984375, output=0.993755553414
			11'd374: out = 32'b00000000000000000111111101000001; // input=1.462890625, output=0.9941838265
			11'd375: out = 32'b00000000000000000111111101001111; // input=1.466796875, output=0.994596929564
			11'd376: out = 32'b00000000000000000111111101011100; // input=1.470703125, output=0.994994856303
			11'd377: out = 32'b00000000000000000111111101101001; // input=1.474609375, output=0.995377600644
			11'd378: out = 32'b00000000000000000111111101110101; // input=1.478515625, output=0.995745156748
			11'd379: out = 32'b00000000000000000111111110000000; // input=1.482421875, output=0.996097519006
			11'd380: out = 32'b00000000000000000111111110001011; // input=1.486328125, output=0.996434682041
			11'd381: out = 32'b00000000000000000111111110010110; // input=1.490234375, output=0.996756640709
			11'd382: out = 32'b00000000000000000111111110100000; // input=1.494140625, output=0.997063390097
			11'd383: out = 32'b00000000000000000111111110101001; // input=1.498046875, output=0.997354925525
			11'd384: out = 32'b00000000000000000111111110110010; // input=1.501953125, output=0.997631242543
			11'd385: out = 32'b00000000000000000111111110111011; // input=1.505859375, output=0.997892336936
			11'd386: out = 32'b00000000000000000111111111000011; // input=1.509765625, output=0.99813820472
			11'd387: out = 32'b00000000000000000111111111001011; // input=1.513671875, output=0.998368842143
			11'd388: out = 32'b00000000000000000111111111010010; // input=1.517578125, output=0.998584245685
			11'd389: out = 32'b00000000000000000111111111011000; // input=1.521484375, output=0.998784412061
			11'd390: out = 32'b00000000000000000111111111011110; // input=1.525390625, output=0.998969338215
			11'd391: out = 32'b00000000000000000111111111100100; // input=1.529296875, output=0.999139021326
			11'd392: out = 32'b00000000000000000111111111101001; // input=1.533203125, output=0.999293458805
			11'd393: out = 32'b00000000000000000111111111101101; // input=1.537109375, output=0.999432648295
			11'd394: out = 32'b00000000000000000111111111110001; // input=1.541015625, output=0.999556587673
			11'd395: out = 32'b00000000000000000111111111110101; // input=1.544921875, output=0.999665275047
			11'd396: out = 32'b00000000000000000111111111111000; // input=1.548828125, output=0.999758708759
			11'd397: out = 32'b00000000000000000111111111111011; // input=1.552734375, output=0.999836887383
			11'd398: out = 32'b00000000000000000111111111111101; // input=1.556640625, output=0.999899809726
			11'd399: out = 32'b00000000000000000111111111111110; // input=1.560546875, output=0.999947474829
			11'd400: out = 32'b00000000000000000111111111111111; // input=1.564453125, output=0.999979881963
			11'd401: out = 32'b00000000000000000111111111111111; // input=1.568359375, output=0.999997030634
			11'd402: out = 32'b00000000000000000111111111111111; // input=1.572265625, output=0.999998920582
			11'd403: out = 32'b00000000000000000111111111111111; // input=1.576171875, output=0.999985551776
			11'd404: out = 32'b00000000000000000111111111111111; // input=1.580078125, output=0.99995692442
			11'd405: out = 32'b00000000000000000111111111111101; // input=1.583984375, output=0.999913038953
			11'd406: out = 32'b00000000000000000111111111111011; // input=1.587890625, output=0.999853896042
			11'd407: out = 32'b00000000000000000111111111111001; // input=1.591796875, output=0.999779496592
			11'd408: out = 32'b00000000000000000111111111110110; // input=1.595703125, output=0.999689841736
			11'd409: out = 32'b00000000000000000111111111110010; // input=1.599609375, output=0.999584932843
			11'd410: out = 32'b00000000000000000111111111101110; // input=1.603515625, output=0.999464771514
			11'd411: out = 32'b00000000000000000111111111101010; // input=1.607421875, output=0.999329359583
			11'd412: out = 32'b00000000000000000111111111100101; // input=1.611328125, output=0.999178699114
			11'd413: out = 32'b00000000000000000111111111100000; // input=1.615234375, output=0.999012792408
			11'd414: out = 32'b00000000000000000111111111011010; // input=1.619140625, output=0.998831641997
			11'd415: out = 32'b00000000000000000111111111010011; // input=1.623046875, output=0.998635250643
			11'd416: out = 32'b00000000000000000111111111001100; // input=1.626953125, output=0.998423621343
			11'd417: out = 32'b00000000000000000111111111000101; // input=1.630859375, output=0.998196757328
			11'd418: out = 32'b00000000000000000111111110111101; // input=1.634765625, output=0.997954662059
			11'd419: out = 32'b00000000000000000111111110110101; // input=1.638671875, output=0.997697339229
			11'd420: out = 32'b00000000000000000111111110101100; // input=1.642578125, output=0.997424792765
			11'd421: out = 32'b00000000000000000111111110100010; // input=1.646484375, output=0.997137026826
			11'd422: out = 32'b00000000000000000111111110011000; // input=1.650390625, output=0.996834045803
			11'd423: out = 32'b00000000000000000111111110001110; // input=1.654296875, output=0.996515854318
			11'd424: out = 32'b00000000000000000111111110000011; // input=1.658203125, output=0.996182457228
			11'd425: out = 32'b00000000000000000111111101110111; // input=1.662109375, output=0.995833859619
			11'd426: out = 32'b00000000000000000111111101101100; // input=1.666015625, output=0.995470066811
			11'd427: out = 32'b00000000000000000111111101011111; // input=1.669921875, output=0.995091084354
			11'd428: out = 32'b00000000000000000111111101010010; // input=1.673828125, output=0.994696918032
			11'd429: out = 32'b00000000000000000111111101000101; // input=1.677734375, output=0.994287573858
			11'd430: out = 32'b00000000000000000111111100110111; // input=1.681640625, output=0.99386305808
			11'd431: out = 32'b00000000000000000111111100101000; // input=1.685546875, output=0.993423377174
			11'd432: out = 32'b00000000000000000111111100011010; // input=1.689453125, output=0.992968537849
			11'd433: out = 32'b00000000000000000111111100001010; // input=1.693359375, output=0.992498547046
			11'd434: out = 32'b00000000000000000111111011111010; // input=1.697265625, output=0.992013411937
			11'd435: out = 32'b00000000000000000111111011101010; // input=1.701171875, output=0.991513139923
			11'd436: out = 32'b00000000000000000111111011011001; // input=1.705078125, output=0.990997738639
			11'd437: out = 32'b00000000000000000111111011001000; // input=1.708984375, output=0.990467215948
			11'd438: out = 32'b00000000000000000111111010110110; // input=1.712890625, output=0.989921579947
			11'd439: out = 32'b00000000000000000111111010100011; // input=1.716796875, output=0.98936083896
			11'd440: out = 32'b00000000000000000111111010010001; // input=1.720703125, output=0.988785001544
			11'd441: out = 32'b00000000000000000111111001111101; // input=1.724609375, output=0.988194076485
			11'd442: out = 32'b00000000000000000111111001101001; // input=1.728515625, output=0.9875880728
			11'd443: out = 32'b00000000000000000111111001010101; // input=1.732421875, output=0.986966999737
			11'd444: out = 32'b00000000000000000111111001000000; // input=1.736328125, output=0.986330866772
			11'd445: out = 32'b00000000000000000111111000101011; // input=1.740234375, output=0.98567968361
			11'd446: out = 32'b00000000000000000111111000010101; // input=1.744140625, output=0.98501346019
			11'd447: out = 32'b00000000000000000111110111111111; // input=1.748046875, output=0.984332206676
			11'd448: out = 32'b00000000000000000111110111101000; // input=1.751953125, output=0.983635933464
			11'd449: out = 32'b00000000000000000111110111010000; // input=1.755859375, output=0.982924651178
			11'd450: out = 32'b00000000000000000111110110111001; // input=1.759765625, output=0.982198370671
			11'd451: out = 32'b00000000000000000111110110100000; // input=1.763671875, output=0.981457103025
			11'd452: out = 32'b00000000000000000111110110001000; // input=1.767578125, output=0.980700859551
			11'd453: out = 32'b00000000000000000111110101101110; // input=1.771484375, output=0.979929651789
			11'd454: out = 32'b00000000000000000111110101010101; // input=1.775390625, output=0.979143491506
			11'd455: out = 32'b00000000000000000111110100111010; // input=1.779296875, output=0.978342390698
			11'd456: out = 32'b00000000000000000111110100100000; // input=1.783203125, output=0.977526361588
			11'd457: out = 32'b00000000000000000111110100000100; // input=1.787109375, output=0.976695416629
			11'd458: out = 32'b00000000000000000111110011101001; // input=1.791015625, output=0.9758495685
			11'd459: out = 32'b00000000000000000111110011001100; // input=1.794921875, output=0.974988830107
			11'd460: out = 32'b00000000000000000111110010110000; // input=1.798828125, output=0.974113214584
			11'd461: out = 32'b00000000000000000111110010010011; // input=1.802734375, output=0.973222735292
			11'd462: out = 32'b00000000000000000111110001110101; // input=1.806640625, output=0.972317405818
			11'd463: out = 32'b00000000000000000111110001010111; // input=1.810546875, output=0.971397239977
			11'd464: out = 32'b00000000000000000111110000111000; // input=1.814453125, output=0.970462251809
			11'd465: out = 32'b00000000000000000111110000011001; // input=1.818359375, output=0.969512455581
			11'd466: out = 32'b00000000000000000111101111111001; // input=1.822265625, output=0.968547865786
			11'd467: out = 32'b00000000000000000111101111011001; // input=1.826171875, output=0.967568497142
			11'd468: out = 32'b00000000000000000111101110111001; // input=1.830078125, output=0.966574364594
			11'd469: out = 32'b00000000000000000111101110011000; // input=1.833984375, output=0.96556548331
			11'd470: out = 32'b00000000000000000111101101110110; // input=1.837890625, output=0.964541868684
			11'd471: out = 32'b00000000000000000111101101010100; // input=1.841796875, output=0.963503536336
			11'd472: out = 32'b00000000000000000111101100110010; // input=1.845703125, output=0.96245050211
			11'd473: out = 32'b00000000000000000111101100001111; // input=1.849609375, output=0.961382782073
			11'd474: out = 32'b00000000000000000111101011101011; // input=1.853515625, output=0.960300392518
			11'd475: out = 32'b00000000000000000111101011000111; // input=1.857421875, output=0.95920334996
			11'd476: out = 32'b00000000000000000111101010100011; // input=1.861328125, output=0.95809167114
			11'd477: out = 32'b00000000000000000111101001111110; // input=1.865234375, output=0.956965373019
			11'd478: out = 32'b00000000000000000111101001011000; // input=1.869140625, output=0.955824472784
			11'd479: out = 32'b00000000000000000111101000110011; // input=1.873046875, output=0.954668987843
			11'd480: out = 32'b00000000000000000111101000001100; // input=1.876953125, output=0.953498935829
			11'd481: out = 32'b00000000000000000111100111100101; // input=1.880859375, output=0.952314334593
			11'd482: out = 32'b00000000000000000111100110111110; // input=1.884765625, output=0.951115202213
			11'd483: out = 32'b00000000000000000111100110010110; // input=1.888671875, output=0.949901556985
			11'd484: out = 32'b00000000000000000111100101101110; // input=1.892578125, output=0.948673417428
			11'd485: out = 32'b00000000000000000111100101000101; // input=1.896484375, output=0.947430802281
			11'd486: out = 32'b00000000000000000111100100011100; // input=1.900390625, output=0.946173730507
			11'd487: out = 32'b00000000000000000111100011110011; // input=1.904296875, output=0.944902221285
			11'd488: out = 32'b00000000000000000111100011001000; // input=1.908203125, output=0.943616294018
			11'd489: out = 32'b00000000000000000111100010011110; // input=1.912109375, output=0.942315968327
			11'd490: out = 32'b00000000000000000111100001110011; // input=1.916015625, output=0.941001264054
			11'd491: out = 32'b00000000000000000111100001000111; // input=1.919921875, output=0.939672201259
			11'd492: out = 32'b00000000000000000111100000011011; // input=1.923828125, output=0.938328800223
			11'd493: out = 32'b00000000000000000111011111101111; // input=1.927734375, output=0.936971081444
			11'd494: out = 32'b00000000000000000111011111000010; // input=1.931640625, output=0.935599065638
			11'd495: out = 32'b00000000000000000111011110010100; // input=1.935546875, output=0.934212773742
			11'd496: out = 32'b00000000000000000111011101100110; // input=1.939453125, output=0.932812226909
			11'd497: out = 32'b00000000000000000111011100111000; // input=1.943359375, output=0.931397446509
			11'd498: out = 32'b00000000000000000111011100001001; // input=1.947265625, output=0.929968454129
			11'd499: out = 32'b00000000000000000111011011011010; // input=1.951171875, output=0.928525271575
			11'd500: out = 32'b00000000000000000111011010101010; // input=1.955078125, output=0.927067920868
			11'd501: out = 32'b00000000000000000111011001111010; // input=1.958984375, output=0.925596424245
			11'd502: out = 32'b00000000000000000111011001001001; // input=1.962890625, output=0.92411080416
			11'd503: out = 32'b00000000000000000111011000011000; // input=1.966796875, output=0.92261108328
			11'd504: out = 32'b00000000000000000111010111100111; // input=1.970703125, output=0.921097284491
			11'd505: out = 32'b00000000000000000111010110110100; // input=1.974609375, output=0.91956943089
			11'd506: out = 32'b00000000000000000111010110000010; // input=1.978515625, output=0.918027545791
			11'd507: out = 32'b00000000000000000111010101001111; // input=1.982421875, output=0.916471652721
			11'd508: out = 32'b00000000000000000111010100011100; // input=1.986328125, output=0.914901775422
			11'd509: out = 32'b00000000000000000111010011101000; // input=1.990234375, output=0.913317937847
			11'd510: out = 32'b00000000000000000111010010110011; // input=1.994140625, output=0.911720164164
			11'd511: out = 32'b00000000000000000111010001111110; // input=1.998046875, output=0.910108478752
			11'd512: out = 32'b00000000000000000111010001001001; // input=2.001953125, output=0.908482906206
			11'd513: out = 32'b00000000000000000111010000010011; // input=2.005859375, output=0.906843471327
			11'd514: out = 32'b00000000000000000111001111011101; // input=2.009765625, output=0.905190199134
			11'd515: out = 32'b00000000000000000111001110100111; // input=2.013671875, output=0.903523114851
			11'd516: out = 32'b00000000000000000111001101110000; // input=2.017578125, output=0.901842243918
			11'd517: out = 32'b00000000000000000111001100111000; // input=2.021484375, output=0.900147611981
			11'd518: out = 32'b00000000000000000111001100000000; // input=2.025390625, output=0.898439244899
			11'd519: out = 32'b00000000000000000111001011001000; // input=2.029296875, output=0.89671716874
			11'd520: out = 32'b00000000000000000111001010001111; // input=2.033203125, output=0.89498140978
			11'd521: out = 32'b00000000000000000111001001010101; // input=2.037109375, output=0.893231994505
			11'd522: out = 32'b00000000000000000111001000011100; // input=2.041015625, output=0.891468949608
			11'd523: out = 32'b00000000000000000111000111100001; // input=2.044921875, output=0.889692301992
			11'd524: out = 32'b00000000000000000111000110100111; // input=2.048828125, output=0.887902078767
			11'd525: out = 32'b00000000000000000111000101101100; // input=2.052734375, output=0.886098307248
			11'd526: out = 32'b00000000000000000111000100110000; // input=2.056640625, output=0.884281014959
			11'd527: out = 32'b00000000000000000111000011110100; // input=2.060546875, output=0.882450229629
			11'd528: out = 32'b00000000000000000111000010111000; // input=2.064453125, output=0.880605979195
			11'd529: out = 32'b00000000000000000111000001111011; // input=2.068359375, output=0.878748291797
			11'd530: out = 32'b00000000000000000111000000111110; // input=2.072265625, output=0.876877195782
			11'd531: out = 32'b00000000000000000111000000000000; // input=2.076171875, output=0.874992719699
			11'd532: out = 32'b00000000000000000110111111000010; // input=2.080078125, output=0.873094892304
			11'd533: out = 32'b00000000000000000110111110000011; // input=2.083984375, output=0.871183742555
			11'd534: out = 32'b00000000000000000110111101000100; // input=2.087890625, output=0.869259299614
			11'd535: out = 32'b00000000000000000110111100000100; // input=2.091796875, output=0.867321592845
			11'd536: out = 32'b00000000000000000110111011000100; // input=2.095703125, output=0.865370651816
			11'd537: out = 32'b00000000000000000110111010000100; // input=2.099609375, output=0.863406506296
			11'd538: out = 32'b00000000000000000110111001000011; // input=2.103515625, output=0.861429186254
			11'd539: out = 32'b00000000000000000110111000000010; // input=2.107421875, output=0.859438721864
			11'd540: out = 32'b00000000000000000110110111000000; // input=2.111328125, output=0.857435143495
			11'd541: out = 32'b00000000000000000110110101111110; // input=2.115234375, output=0.855418481721
			11'd542: out = 32'b00000000000000000110110100111100; // input=2.119140625, output=0.853388767314
			11'd543: out = 32'b00000000000000000110110011111001; // input=2.123046875, output=0.851346031244
			11'd544: out = 32'b00000000000000000110110010110110; // input=2.126953125, output=0.849290304681
			11'd545: out = 32'b00000000000000000110110001110010; // input=2.130859375, output=0.847221618993
			11'd546: out = 32'b00000000000000000110110000101110; // input=2.134765625, output=0.845140005746
			11'd547: out = 32'b00000000000000000110101111101001; // input=2.138671875, output=0.843045496701
			11'd548: out = 32'b00000000000000000110101110100100; // input=2.142578125, output=0.84093812382
			11'd549: out = 32'b00000000000000000110101101011110; // input=2.146484375, output=0.838817919257
			11'd550: out = 32'b00000000000000000110101100011000; // input=2.150390625, output=0.836684915366
			11'd551: out = 32'b00000000000000000110101011010010; // input=2.154296875, output=0.834539144691
			11'd552: out = 32'b00000000000000000110101010001011; // input=2.158203125, output=0.832380639976
			11'd553: out = 32'b00000000000000000110101001000100; // input=2.162109375, output=0.830209434157
			11'd554: out = 32'b00000000000000000110100111111101; // input=2.166015625, output=0.828025560363
			11'd555: out = 32'b00000000000000000110100110110101; // input=2.169921875, output=0.825829051918
			11'd556: out = 32'b00000000000000000110100101101100; // input=2.173828125, output=0.823619942338
			11'd557: out = 32'b00000000000000000110100100100100; // input=2.177734375, output=0.82139826533
			11'd558: out = 32'b00000000000000000110100011011010; // input=2.181640625, output=0.819164054796
			11'd559: out = 32'b00000000000000000110100010010001; // input=2.185546875, output=0.816917344826
			11'd560: out = 32'b00000000000000000110100001000111; // input=2.189453125, output=0.814658169702
			11'd561: out = 32'b00000000000000000110011111111100; // input=2.193359375, output=0.812386563897
			11'd562: out = 32'b00000000000000000110011110110001; // input=2.197265625, output=0.810102562073
			11'd563: out = 32'b00000000000000000110011101100110; // input=2.201171875, output=0.80780619908
			11'd564: out = 32'b00000000000000000110011100011011; // input=2.205078125, output=0.805497509959
			11'd565: out = 32'b00000000000000000110011011001110; // input=2.208984375, output=0.803176529936
			11'd566: out = 32'b00000000000000000110011010000010; // input=2.212890625, output=0.800843294428
			11'd567: out = 32'b00000000000000000110011000110101; // input=2.216796875, output=0.798497839037
			11'd568: out = 32'b00000000000000000110010111101000; // input=2.220703125, output=0.796140199551
			11'd569: out = 32'b00000000000000000110010110011010; // input=2.224609375, output=0.793770411945
			11'd570: out = 32'b00000000000000000110010101001100; // input=2.228515625, output=0.791388512379
			11'd571: out = 32'b00000000000000000110010011111110; // input=2.232421875, output=0.788994537198
			11'd572: out = 32'b00000000000000000110010010101111; // input=2.236328125, output=0.786588522931
			11'd573: out = 32'b00000000000000000110010001100000; // input=2.240234375, output=0.784170506291
			11'd574: out = 32'b00000000000000000110010000010000; // input=2.244140625, output=0.781740524174
			11'd575: out = 32'b00000000000000000110001111000000; // input=2.248046875, output=0.779298613658
			11'd576: out = 32'b00000000000000000110001101110000; // input=2.251953125, output=0.776844812005
			11'd577: out = 32'b00000000000000000110001100011111; // input=2.255859375, output=0.774379156655
			11'd578: out = 32'b00000000000000000110001011001110; // input=2.259765625, output=0.771901685232
			11'd579: out = 32'b00000000000000000110001001111100; // input=2.263671875, output=0.769412435539
			11'd580: out = 32'b00000000000000000110001000101010; // input=2.267578125, output=0.766911445559
			11'd581: out = 32'b00000000000000000110000111011000; // input=2.271484375, output=0.764398753454
			11'd582: out = 32'b00000000000000000110000110000101; // input=2.275390625, output=0.761874397564
			11'd583: out = 32'b00000000000000000110000100110010; // input=2.279296875, output=0.759338416409
			11'd584: out = 32'b00000000000000000110000011011111; // input=2.283203125, output=0.756790848683
			11'd585: out = 32'b00000000000000000110000010001011; // input=2.287109375, output=0.75423173326
			11'd586: out = 32'b00000000000000000110000000110110; // input=2.291015625, output=0.751661109189
			11'd587: out = 32'b00000000000000000101111111100010; // input=2.294921875, output=0.749079015694
			11'd588: out = 32'b00000000000000000101111110001101; // input=2.298828125, output=0.746485492175
			11'd589: out = 32'b00000000000000000101111100110111; // input=2.302734375, output=0.743880578206
			11'd590: out = 32'b00000000000000000101111011100010; // input=2.306640625, output=0.741264313535
			11'd591: out = 32'b00000000000000000101111010001100; // input=2.310546875, output=0.738636738082
			11'd592: out = 32'b00000000000000000101111000110101; // input=2.314453125, output=0.735997891941
			11'd593: out = 32'b00000000000000000101110111011110; // input=2.318359375, output=0.733347815378
			11'd594: out = 32'b00000000000000000101110110000111; // input=2.322265625, output=0.730686548829
			11'd595: out = 32'b00000000000000000101110100110000; // input=2.326171875, output=0.728014132903
			11'd596: out = 32'b00000000000000000101110011011000; // input=2.330078125, output=0.725330608377
			11'd597: out = 32'b00000000000000000101110001111111; // input=2.333984375, output=0.722636016198
			11'd598: out = 32'b00000000000000000101110000100111; // input=2.337890625, output=0.719930397482
			11'd599: out = 32'b00000000000000000101101111001110; // input=2.341796875, output=0.717213793515
			11'd600: out = 32'b00000000000000000101101101110100; // input=2.345703125, output=0.714486245747
			11'd601: out = 32'b00000000000000000101101100011011; // input=2.349609375, output=0.711747795798
			11'd602: out = 32'b00000000000000000101101011000000; // input=2.353515625, output=0.708998485454
			11'd603: out = 32'b00000000000000000101101001100110; // input=2.357421875, output=0.706238356665
			11'd604: out = 32'b00000000000000000101101000001011; // input=2.361328125, output=0.703467451548
			11'd605: out = 32'b00000000000000000101100110110000; // input=2.365234375, output=0.700685812383
			11'd606: out = 32'b00000000000000000101100101010101; // input=2.369140625, output=0.697893481614
			11'd607: out = 32'b00000000000000000101100011111001; // input=2.373046875, output=0.69509050185
			11'd608: out = 32'b00000000000000000101100010011101; // input=2.376953125, output=0.692276915859
			11'd609: out = 32'b00000000000000000101100001000000; // input=2.380859375, output=0.689452766575
			11'd610: out = 32'b00000000000000000101011111100011; // input=2.384765625, output=0.68661809709
			11'd611: out = 32'b00000000000000000101011110000110; // input=2.388671875, output=0.683772950657
			11'd612: out = 32'b00000000000000000101011100101000; // input=2.392578125, output=0.680917370691
			11'd613: out = 32'b00000000000000000101011011001010; // input=2.396484375, output=0.678051400763
			11'd614: out = 32'b00000000000000000101011001101100; // input=2.400390625, output=0.675175084605
			11'd615: out = 32'b00000000000000000101011000001110; // input=2.404296875, output=0.672288466105
			11'd616: out = 32'b00000000000000000101010110101111; // input=2.408203125, output=0.669391589311
			11'd617: out = 32'b00000000000000000101010101001111; // input=2.412109375, output=0.666484498425
			11'd618: out = 32'b00000000000000000101010011110000; // input=2.416015625, output=0.663567237806
			11'd619: out = 32'b00000000000000000101010010010000; // input=2.419921875, output=0.660639851967
			11'd620: out = 32'b00000000000000000101010000110000; // input=2.423828125, output=0.657702385576
			11'd621: out = 32'b00000000000000000101001111001111; // input=2.427734375, output=0.654754883457
			11'd622: out = 32'b00000000000000000101001101101110; // input=2.431640625, output=0.651797390583
			11'd623: out = 32'b00000000000000000101001100001101; // input=2.435546875, output=0.648829952083
			11'd624: out = 32'b00000000000000000101001010101011; // input=2.439453125, output=0.645852613236
			11'd625: out = 32'b00000000000000000101001001001001; // input=2.443359375, output=0.642865419473
			11'd626: out = 32'b00000000000000000101000111100111; // input=2.447265625, output=0.639868416375
			11'd627: out = 32'b00000000000000000101000110000101; // input=2.451171875, output=0.636861649672
			11'd628: out = 32'b00000000000000000101000100100010; // input=2.455078125, output=0.633845165244
			11'd629: out = 32'b00000000000000000101000010111111; // input=2.458984375, output=0.630819009118
			11'd630: out = 32'b00000000000000000101000001011011; // input=2.462890625, output=0.62778322747
			11'd631: out = 32'b00000000000000000100111111110111; // input=2.466796875, output=0.624737866623
			11'd632: out = 32'b00000000000000000100111110010011; // input=2.470703125, output=0.621682973045
			11'd633: out = 32'b00000000000000000100111100101111; // input=2.474609375, output=0.618618593349
			11'd634: out = 32'b00000000000000000100111011001010; // input=2.478515625, output=0.615544774295
			11'd635: out = 32'b00000000000000000100111001100101; // input=2.482421875, output=0.612461562784
			11'd636: out = 32'b00000000000000000100111000000000; // input=2.486328125, output=0.609369005864
			11'd637: out = 32'b00000000000000000100110110011010; // input=2.490234375, output=0.606267150722
			11'd638: out = 32'b00000000000000000100110100110100; // input=2.494140625, output=0.60315604469
			11'd639: out = 32'b00000000000000000100110011001110; // input=2.498046875, output=0.600035735239
			11'd640: out = 32'b00000000000000000100110001100111; // input=2.501953125, output=0.59690626998
			11'd641: out = 32'b00000000000000000100110000000001; // input=2.505859375, output=0.593767696666
			11'd642: out = 32'b00000000000000000100101110011001; // input=2.509765625, output=0.590620063188
			11'd643: out = 32'b00000000000000000100101100110010; // input=2.513671875, output=0.587463417574
			11'd644: out = 32'b00000000000000000100101011001010; // input=2.517578125, output=0.584297807991
			11'd645: out = 32'b00000000000000000100101001100010; // input=2.521484375, output=0.581123282743
			11'd646: out = 32'b00000000000000000100100111111010; // input=2.525390625, output=0.577939890268
			11'd647: out = 32'b00000000000000000100100110010001; // input=2.529296875, output=0.574747679141
			11'd648: out = 32'b00000000000000000100100100101000; // input=2.533203125, output=0.571546698072
			11'd649: out = 32'b00000000000000000100100010111111; // input=2.537109375, output=0.568336995904
			11'd650: out = 32'b00000000000000000100100001010110; // input=2.541015625, output=0.565118621612
			11'd651: out = 32'b00000000000000000100011111101100; // input=2.544921875, output=0.561891624306
			11'd652: out = 32'b00000000000000000100011110000010; // input=2.548828125, output=0.558656053224
			11'd653: out = 32'b00000000000000000100011100011000; // input=2.552734375, output=0.555411957739
			11'd654: out = 32'b00000000000000000100011010101101; // input=2.556640625, output=0.55215938735
			11'd655: out = 32'b00000000000000000100011001000010; // input=2.560546875, output=0.548898391689
			11'd656: out = 32'b00000000000000000100010111010111; // input=2.564453125, output=0.545629020513
			11'd657: out = 32'b00000000000000000100010101101100; // input=2.568359375, output=0.54235132371
			11'd658: out = 32'b00000000000000000100010100000000; // input=2.572265625, output=0.539065351293
			11'd659: out = 32'b00000000000000000100010010010100; // input=2.576171875, output=0.535771153402
			11'd660: out = 32'b00000000000000000100010000101000; // input=2.580078125, output=0.532468780302
			11'd661: out = 32'b00000000000000000100001110111011; // input=2.583984375, output=0.529158282384
			11'd662: out = 32'b00000000000000000100001101001111; // input=2.587890625, output=0.525839710162
			11'd663: out = 32'b00000000000000000100001011100010; // input=2.591796875, output=0.522513114272
			11'd664: out = 32'b00000000000000000100001001110100; // input=2.595703125, output=0.519178545475
			11'd665: out = 32'b00000000000000000100001000000111; // input=2.599609375, output=0.515836054653
			11'd666: out = 32'b00000000000000000100000110011001; // input=2.603515625, output=0.512485692806
			11'd667: out = 32'b00000000000000000100000100101011; // input=2.607421875, output=0.509127511059
			11'd668: out = 32'b00000000000000000100000010111101; // input=2.611328125, output=0.505761560652
			11'd669: out = 32'b00000000000000000100000001001110; // input=2.615234375, output=0.502387892946
			11'd670: out = 32'b00000000000000000011111111011111; // input=2.619140625, output=0.499006559419
			11'd671: out = 32'b00000000000000000011111101110000; // input=2.623046875, output=0.495617611666
			11'd672: out = 32'b00000000000000000011111100000001; // input=2.626953125, output=0.492221101398
			11'd673: out = 32'b00000000000000000011111010010010; // input=2.630859375, output=0.488817080442
			11'd674: out = 32'b00000000000000000011111000100010; // input=2.634765625, output=0.485405600738
			11'd675: out = 32'b00000000000000000011110110110010; // input=2.638671875, output=0.481986714342
			11'd676: out = 32'b00000000000000000011110101000001; // input=2.642578125, output=0.478560473421
			11'd677: out = 32'b00000000000000000011110011010001; // input=2.646484375, output=0.475126930257
			11'd678: out = 32'b00000000000000000011110001100000; // input=2.650390625, output=0.47168613724
			11'd679: out = 32'b00000000000000000011101111101111; // input=2.654296875, output=0.468238146873
			11'd680: out = 32'b00000000000000000011101101111110; // input=2.658203125, output=0.464783011769
			11'd681: out = 32'b00000000000000000011101100001101; // input=2.662109375, output=0.461320784647
			11'd682: out = 32'b00000000000000000011101010011011; // input=2.666015625, output=0.457851518337
			11'd683: out = 32'b00000000000000000011101000101001; // input=2.669921875, output=0.454375265777
			11'd684: out = 32'b00000000000000000011100110110111; // input=2.673828125, output=0.450892080009
			11'd685: out = 32'b00000000000000000011100101000100; // input=2.677734375, output=0.447402014183
			11'd686: out = 32'b00000000000000000011100011010010; // input=2.681640625, output=0.443905121553
			11'd687: out = 32'b00000000000000000011100001011111; // input=2.685546875, output=0.440401455476
			11'd688: out = 32'b00000000000000000011011111101100; // input=2.689453125, output=0.436891069416
			11'd689: out = 32'b00000000000000000011011101111001; // input=2.693359375, output=0.433374016935
			11'd690: out = 32'b00000000000000000011011100000101; // input=2.697265625, output=0.429850351699
			11'd691: out = 32'b00000000000000000011011010010010; // input=2.701171875, output=0.426320127476
			11'd692: out = 32'b00000000000000000011011000011110; // input=2.705078125, output=0.422783398133
			11'd693: out = 32'b00000000000000000011010110101010; // input=2.708984375, output=0.419240217635
			11'd694: out = 32'b00000000000000000011010100110101; // input=2.712890625, output=0.415690640047
			11'd695: out = 32'b00000000000000000011010011000001; // input=2.716796875, output=0.412134719532
			11'd696: out = 32'b00000000000000000011010001001100; // input=2.720703125, output=0.408572510347
			11'd697: out = 32'b00000000000000000011001111010111; // input=2.724609375, output=0.405004066849
			11'd698: out = 32'b00000000000000000011001101100010; // input=2.728515625, output=0.401429443487
			11'd699: out = 32'b00000000000000000011001011101101; // input=2.732421875, output=0.397848694806
			11'd700: out = 32'b00000000000000000011001001110111; // input=2.736328125, output=0.394261875443
			11'd701: out = 32'b00000000000000000011001000000001; // input=2.740234375, output=0.390669040129
			11'd702: out = 32'b00000000000000000011000110001100; // input=2.744140625, output=0.387070243686
			11'd703: out = 32'b00000000000000000011000100010101; // input=2.748046875, output=0.383465541027
			11'd704: out = 32'b00000000000000000011000010011111; // input=2.751953125, output=0.379854987156
			11'd705: out = 32'b00000000000000000011000000101001; // input=2.755859375, output=0.376238637166
			11'd706: out = 32'b00000000000000000010111110110010; // input=2.759765625, output=0.372616546236
			11'd707: out = 32'b00000000000000000010111100111011; // input=2.763671875, output=0.368988769637
			11'd708: out = 32'b00000000000000000010111011000100; // input=2.767578125, output=0.365355362723
			11'd709: out = 32'b00000000000000000010111001001101; // input=2.771484375, output=0.361716380935
			11'd710: out = 32'b00000000000000000010110111010101; // input=2.775390625, output=0.358071879801
			11'd711: out = 32'b00000000000000000010110101011110; // input=2.779296875, output=0.35442191493
			11'd712: out = 32'b00000000000000000010110011100110; // input=2.783203125, output=0.350766542017
			11'd713: out = 32'b00000000000000000010110001101110; // input=2.787109375, output=0.347105816838
			11'd714: out = 32'b00000000000000000010101111110110; // input=2.791015625, output=0.343439795251
			11'd715: out = 32'b00000000000000000010101101111110; // input=2.794921875, output=0.339768533196
			11'd716: out = 32'b00000000000000000010101100000101; // input=2.798828125, output=0.336092086691
			11'd717: out = 32'b00000000000000000010101010001100; // input=2.802734375, output=0.332410511834
			11'd718: out = 32'b00000000000000000010101000010100; // input=2.806640625, output=0.328723864801
			11'd719: out = 32'b00000000000000000010100110011011; // input=2.810546875, output=0.325032201847
			11'd720: out = 32'b00000000000000000010100100100010; // input=2.814453125, output=0.321335579302
			11'd721: out = 32'b00000000000000000010100010101000; // input=2.818359375, output=0.31763405357
			11'd722: out = 32'b00000000000000000010100000101111; // input=2.822265625, output=0.313927681134
			11'd723: out = 32'b00000000000000000010011110110101; // input=2.826171875, output=0.310216518548
			11'd724: out = 32'b00000000000000000010011100111011; // input=2.830078125, output=0.306500622439
			11'd725: out = 32'b00000000000000000010011011000001; // input=2.833984375, output=0.302780049508
			11'd726: out = 32'b00000000000000000010011001000111; // input=2.837890625, output=0.299054856526
			11'd727: out = 32'b00000000000000000010010111001101; // input=2.841796875, output=0.295325100335
			11'd728: out = 32'b00000000000000000010010101010011; // input=2.845703125, output=0.291590837846
			11'd729: out = 32'b00000000000000000010010011011000; // input=2.849609375, output=0.28785212604
			11'd730: out = 32'b00000000000000000010010001011110; // input=2.853515625, output=0.284109021964
			11'd731: out = 32'b00000000000000000010001111100011; // input=2.857421875, output=0.280361582734
			11'd732: out = 32'b00000000000000000010001101101000; // input=2.861328125, output=0.276609865532
			11'd733: out = 32'b00000000000000000010001011101101; // input=2.865234375, output=0.272853927603
			11'd734: out = 32'b00000000000000000010001001110010; // input=2.869140625, output=0.269093826259
			11'd735: out = 32'b00000000000000000010000111110110; // input=2.873046875, output=0.265329618874
			11'd736: out = 32'b00000000000000000010000101111011; // input=2.876953125, output=0.261561362886
			11'd737: out = 32'b00000000000000000010000011111111; // input=2.880859375, output=0.257789115793
			11'd738: out = 32'b00000000000000000010000010000011; // input=2.884765625, output=0.254012935156
			11'd739: out = 32'b00000000000000000010000000001000; // input=2.888671875, output=0.250232878593
			11'd740: out = 32'b00000000000000000001111110001100; // input=2.892578125, output=0.246449003785
			11'd741: out = 32'b00000000000000000001111100010000; // input=2.896484375, output=0.242661368468
			11'd742: out = 32'b00000000000000000001111010010011; // input=2.900390625, output=0.238870030437
			11'd743: out = 32'b00000000000000000001111000010111; // input=2.904296875, output=0.235075047543
			11'd744: out = 32'b00000000000000000001110110011010; // input=2.908203125, output=0.231276477694
			11'd745: out = 32'b00000000000000000001110100011110; // input=2.912109375, output=0.22747437885
			11'd746: out = 32'b00000000000000000001110010100001; // input=2.916015625, output=0.223668809027
			11'd747: out = 32'b00000000000000000001110000100100; // input=2.919921875, output=0.219859826292
			11'd748: out = 32'b00000000000000000001101110100111; // input=2.923828125, output=0.216047488768
			11'd749: out = 32'b00000000000000000001101100101010; // input=2.927734375, output=0.212231854624
			11'd750: out = 32'b00000000000000000001101010101101; // input=2.931640625, output=0.208412982084
			11'd751: out = 32'b00000000000000000001101000110000; // input=2.935546875, output=0.204590929418
			11'd752: out = 32'b00000000000000000001100110110011; // input=2.939453125, output=0.200765754946
			11'd753: out = 32'b00000000000000000001100100110101; // input=2.943359375, output=0.196937517036
			11'd754: out = 32'b00000000000000000001100010111000; // input=2.947265625, output=0.193106274101
			11'd755: out = 32'b00000000000000000001100000111010; // input=2.951171875, output=0.189272084602
			11'd756: out = 32'b00000000000000000001011110111100; // input=2.955078125, output=0.185435007044
			11'd757: out = 32'b00000000000000000001011100111111; // input=2.958984375, output=0.181595099977
			11'd758: out = 32'b00000000000000000001011011000001; // input=2.962890625, output=0.177752421991
			11'd759: out = 32'b00000000000000000001011001000011; // input=2.966796875, output=0.173907031722
			11'd760: out = 32'b00000000000000000001010111000100; // input=2.970703125, output=0.170058987846
			11'd761: out = 32'b00000000000000000001010101000110; // input=2.974609375, output=0.166208349078
			11'd762: out = 32'b00000000000000000001010011001000; // input=2.978515625, output=0.162355174176
			11'd763: out = 32'b00000000000000000001010001001010; // input=2.982421875, output=0.158499521934
			11'd764: out = 32'b00000000000000000001001111001011; // input=2.986328125, output=0.154641451184
			11'd765: out = 32'b00000000000000000001001101001101; // input=2.990234375, output=0.150781020795
			11'd766: out = 32'b00000000000000000001001011001110; // input=2.994140625, output=0.146918289674
			11'd767: out = 32'b00000000000000000001001001010000; // input=2.998046875, output=0.14305331676
			11'd768: out = 32'b00000000000000000001000111010001; // input=3.001953125, output=0.139186161029
			11'd769: out = 32'b00000000000000000001000101010010; // input=3.005859375, output=0.135316881489
			11'd770: out = 32'b00000000000000000001000011010011; // input=3.009765625, output=0.131445537179
			11'd771: out = 32'b00000000000000000001000001010100; // input=3.013671875, output=0.127572187172
			11'd772: out = 32'b00000000000000000000111111010101; // input=3.017578125, output=0.12369689057
			11'd773: out = 32'b00000000000000000000111101010110; // input=3.021484375, output=0.119819706506
			11'd774: out = 32'b00000000000000000000111011010111; // input=3.025390625, output=0.115940694141
			11'd775: out = 32'b00000000000000000000111001011000; // input=3.029296875, output=0.112059912663
			11'd776: out = 32'b00000000000000000000110111011001; // input=3.033203125, output=0.108177421289
			11'd777: out = 32'b00000000000000000000110101011001; // input=3.037109375, output=0.10429327926
			11'd778: out = 32'b00000000000000000000110011011010; // input=3.041015625, output=0.100407545845
			11'd779: out = 32'b00000000000000000000110001011011; // input=3.044921875, output=0.0965202803338
			11'd780: out = 32'b00000000000000000000101111011011; // input=3.048828125, output=0.0926315420419
			11'd781: out = 32'b00000000000000000000101101011100; // input=3.052734375, output=0.0887413903066
			11'd782: out = 32'b00000000000000000000101011011100; // input=3.056640625, output=0.0848498844869
			11'd783: out = 32'b00000000000000000000101001011101; // input=3.060546875, output=0.0809570839624
			11'd784: out = 32'b00000000000000000000100111011101; // input=3.064453125, output=0.0770630481324
			11'd785: out = 32'b00000000000000000000100101011110; // input=3.068359375, output=0.0731678364151
			11'd786: out = 32'b00000000000000000000100011011110; // input=3.072265625, output=0.0692715082466
			11'd787: out = 32'b00000000000000000000100001011110; // input=3.076171875, output=0.0653741230801
			11'd788: out = 32'b00000000000000000000011111011110; // input=3.080078125, output=0.061475740385
			11'd789: out = 32'b00000000000000000000011101011111; // input=3.083984375, output=0.0575764196456
			11'd790: out = 32'b00000000000000000000011011011111; // input=3.087890625, output=0.053676220361
			11'd791: out = 32'b00000000000000000000011001011111; // input=3.091796875, output=0.0497752020432
			11'd792: out = 32'b00000000000000000000010111011111; // input=3.095703125, output=0.0458734242172
			11'd793: out = 32'b00000000000000000000010101011111; // input=3.099609375, output=0.0419709464191
			11'd794: out = 32'b00000000000000000000010011011111; // input=3.103515625, output=0.038067828196
			11'd795: out = 32'b00000000000000000000010001011111; // input=3.107421875, output=0.0341641291047
			11'd796: out = 32'b00000000000000000000001111100000; // input=3.111328125, output=0.0302599087108
			11'd797: out = 32'b00000000000000000000001101100000; // input=3.115234375, output=0.0263552265879
			11'd798: out = 32'b00000000000000000000001011100000; // input=3.119140625, output=0.0224501423167
			11'd799: out = 32'b00000000000000000000001001100000; // input=3.123046875, output=0.018544715484
			11'd800: out = 32'b00000000000000000000000111100000; // input=3.126953125, output=0.0146390056817
			11'd801: out = 32'b00000000000000000000000101100000; // input=3.130859375, output=0.0107330725062
			11'd802: out = 32'b00000000000000000000000011100000; // input=3.134765625, output=0.0068269755572
			11'd803: out = 32'b00000000000000000000000001100000; // input=3.138671875, output=0.00292077443696
			11'd804: out = 32'b10000000000000000000000000100000; // input=3.142578125, output=-0.000985471250699
			11'd805: out = 32'b10000000000000000000000010100000; // input=3.146484375, output=-0.00489170190128
			11'd806: out = 32'b10000000000000000000000100100000; // input=3.150390625, output=-0.00879785791051
			11'd807: out = 32'b10000000000000000000000110100000; // input=3.154296875, output=-0.0127038796752
			11'd808: out = 32'b10000000000000000000001000100000; // input=3.158203125, output=-0.0166097075944
			11'd809: out = 32'b10000000000000000000001010100000; // input=3.162109375, output=-0.0205152820699
			11'd810: out = 32'b10000000000000000000001100100000; // input=3.166015625, output=-0.0244205435074
			11'd811: out = 32'b10000000000000000000001110100000; // input=3.169921875, output=-0.0283254323174
			11'd812: out = 32'b10000000000000000000010000100000; // input=3.173828125, output=-0.0322298889162
			11'd813: out = 32'b10000000000000000000010010100000; // input=3.177734375, output=-0.0361338537266
			11'd814: out = 32'b10000000000000000000010100100000; // input=3.181640625, output=-0.0400372671788
			11'd815: out = 32'b10000000000000000000010110100000; // input=3.185546875, output=-0.0439400697116
			11'd816: out = 32'b10000000000000000000011000100000; // input=3.189453125, output=-0.0478422017729
			11'd817: out = 32'b10000000000000000000011010100000; // input=3.193359375, output=-0.0517436038212
			11'd818: out = 32'b10000000000000000000011100011111; // input=3.197265625, output=-0.0556442163256
			11'd819: out = 32'b10000000000000000000011110011111; // input=3.201171875, output=-0.0595439797679
			11'd820: out = 32'b10000000000000000000100000011111; // input=3.205078125, output=-0.0634428346422
			11'd821: out = 32'b10000000000000000000100010011111; // input=3.208984375, output=-0.0673407214569
			11'd822: out = 32'b10000000000000000000100100011110; // input=3.212890625, output=-0.0712375807351
			11'd823: out = 32'b10000000000000000000100110011110; // input=3.216796875, output=-0.0751333530155
			11'd824: out = 32'b10000000000000000000101000011110; // input=3.220703125, output=-0.0790279788533
			11'd825: out = 32'b10000000000000000000101010011101; // input=3.224609375, output=-0.0829213988214
			11'd826: out = 32'b10000000000000000000101100011101; // input=3.228515625, output=-0.086813553511
			11'd827: out = 32'b10000000000000000000101110011100; // input=3.232421875, output=-0.0907043835325
			11'd828: out = 32'b10000000000000000000110000011100; // input=3.236328125, output=-0.0945938295168
			11'd829: out = 32'b10000000000000000000110010011011; // input=3.240234375, output=-0.0984818321156
			11'd830: out = 32'b10000000000000000000110100011010; // input=3.244140625, output=-0.102368332003
			11'd831: out = 32'b10000000000000000000110110011010; // input=3.248046875, output=-0.106253269875
			11'd832: out = 32'b10000000000000000000111000011001; // input=3.251953125, output=-0.110136586453
			11'd833: out = 32'b10000000000000000000111010011000; // input=3.255859375, output=-0.114018222483
			11'd834: out = 32'b10000000000000000000111100010111; // input=3.259765625, output=-0.117898118735
			11'd835: out = 32'b10000000000000000000111110010110; // input=3.263671875, output=-0.121776216006
			11'd836: out = 32'b10000000000000000001000000010101; // input=3.267578125, output=-0.125652455122
			11'd837: out = 32'b10000000000000000001000010010100; // input=3.271484375, output=-0.129526776936
			11'd838: out = 32'b10000000000000000001000100010011; // input=3.275390625, output=-0.133399122331
			11'd839: out = 32'b10000000000000000001000110010010; // input=3.279296875, output=-0.13726943222
			11'd840: out = 32'b10000000000000000001001000010001; // input=3.283203125, output=-0.141137647546
			11'd841: out = 32'b10000000000000000001001010001111; // input=3.287109375, output=-0.145003709285
			11'd842: out = 32'b10000000000000000001001100001110; // input=3.291015625, output=-0.148867558446
			11'd843: out = 32'b10000000000000000001001110001101; // input=3.294921875, output=-0.152729136071
			11'd844: out = 32'b10000000000000000001010000001011; // input=3.298828125, output=-0.156588383237
			11'd845: out = 32'b10000000000000000001010010001001; // input=3.302734375, output=-0.160445241058
			11'd846: out = 32'b10000000000000000001010100001000; // input=3.306640625, output=-0.164299650681
			11'd847: out = 32'b10000000000000000001010110000110; // input=3.310546875, output=-0.168151553294
			11'd848: out = 32'b10000000000000000001011000000100; // input=3.314453125, output=-0.172000890121
			11'd849: out = 32'b10000000000000000001011010000010; // input=3.318359375, output=-0.175847602426
			11'd850: out = 32'b10000000000000000001011100000000; // input=3.322265625, output=-0.179691631513
			11'd851: out = 32'b10000000000000000001011101111110; // input=3.326171875, output=-0.183532918727
			11'd852: out = 32'b10000000000000000001011111111100; // input=3.330078125, output=-0.187371405454
			11'd853: out = 32'b10000000000000000001100001111001; // input=3.333984375, output=-0.191207033124
			11'd854: out = 32'b10000000000000000001100011110111; // input=3.337890625, output=-0.19503974321
			11'd855: out = 32'b10000000000000000001100101110101; // input=3.341796875, output=-0.198869477229
			11'd856: out = 32'b10000000000000000001100111110010; // input=3.345703125, output=-0.202696176745
			11'd857: out = 32'b10000000000000000001101001101111; // input=3.349609375, output=-0.206519783367
			11'd858: out = 32'b10000000000000000001101011101100; // input=3.353515625, output=-0.210340238751
			11'd859: out = 32'b10000000000000000001101101101010; // input=3.357421875, output=-0.214157484602
			11'd860: out = 32'b10000000000000000001101111100110; // input=3.361328125, output=-0.217971462672
			11'd861: out = 32'b10000000000000000001110001100011; // input=3.365234375, output=-0.221782114767
			11'd862: out = 32'b10000000000000000001110011100000; // input=3.369140625, output=-0.225589382739
			11'd863: out = 32'b10000000000000000001110101011101; // input=3.373046875, output=-0.229393208495
			11'd864: out = 32'b10000000000000000001110111011001; // input=3.376953125, output=-0.233193533993
			11'd865: out = 32'b10000000000000000001111001010110; // input=3.380859375, output=-0.236990301245
			11'd866: out = 32'b10000000000000000001111011010010; // input=3.384765625, output=-0.240783452315
			11'd867: out = 32'b10000000000000000001111101001110; // input=3.388671875, output=-0.244572929327
			11'd868: out = 32'b10000000000000000001111111001010; // input=3.392578125, output=-0.248358674457
			11'd869: out = 32'b10000000000000000010000001000110; // input=3.396484375, output=-0.252140629939
			11'd870: out = 32'b10000000000000000010000011000010; // input=3.400390625, output=-0.255918738065
			11'd871: out = 32'b10000000000000000010000100111110; // input=3.404296875, output=-0.259692941186
			11'd872: out = 32'b10000000000000000010000110111001; // input=3.408203125, output=-0.263463181712
			11'd873: out = 32'b10000000000000000010001000110101; // input=3.412109375, output=-0.267229402115
			11'd874: out = 32'b10000000000000000010001010110000; // input=3.416015625, output=-0.270991544925
			11'd875: out = 32'b10000000000000000010001100101011; // input=3.419921875, output=-0.274749552738
			11'd876: out = 32'b10000000000000000010001110100110; // input=3.423828125, output=-0.27850336821
			11'd877: out = 32'b10000000000000000010010000100001; // input=3.427734375, output=-0.282252934064
			11'd878: out = 32'b10000000000000000010010010011100; // input=3.431640625, output=-0.285998193086
			11'd879: out = 32'b10000000000000000010010100010110; // input=3.435546875, output=-0.289739088127
			11'd880: out = 32'b10000000000000000010010110010001; // input=3.439453125, output=-0.293475562106
			11'd881: out = 32'b10000000000000000010011000001011; // input=3.443359375, output=-0.297207558008
			11'd882: out = 32'b10000000000000000010011010000101; // input=3.447265625, output=-0.30093501889
			11'd883: out = 32'b10000000000000000010011011111111; // input=3.451171875, output=-0.304657887873
			11'd884: out = 32'b10000000000000000010011101111001; // input=3.455078125, output=-0.308376108151
			11'd885: out = 32'b10000000000000000010011111110011; // input=3.458984375, output=-0.31208962299
			11'd886: out = 32'b10000000000000000010100001101100; // input=3.462890625, output=-0.315798375725
			11'd887: out = 32'b10000000000000000010100011100101; // input=3.466796875, output=-0.319502309765
			11'd888: out = 32'b10000000000000000010100101011111; // input=3.470703125, output=-0.323201368593
			11'd889: out = 32'b10000000000000000010100111011000; // input=3.474609375, output=-0.326895495766
			11'd890: out = 32'b10000000000000000010101001010001; // input=3.478515625, output=-0.330584634915
			11'd891: out = 32'b10000000000000000010101011001001; // input=3.482421875, output=-0.33426872975
			11'd892: out = 32'b10000000000000000010101101000010; // input=3.486328125, output=-0.337947724056
			11'd893: out = 32'b10000000000000000010101110111010; // input=3.490234375, output=-0.341621561694
			11'd894: out = 32'b10000000000000000010110000110010; // input=3.494140625, output=-0.345290186609
			11'd895: out = 32'b10000000000000000010110010101011; // input=3.498046875, output=-0.348953542819
			11'd896: out = 32'b10000000000000000010110100100010; // input=3.501953125, output=-0.352611574428
			11'd897: out = 32'b10000000000000000010110110011010; // input=3.505859375, output=-0.356264225619
			11'd898: out = 32'b10000000000000000010111000010010; // input=3.509765625, output=-0.359911440655
			11'd899: out = 32'b10000000000000000010111010001001; // input=3.513671875, output=-0.363553163886
			11'd900: out = 32'b10000000000000000010111100000000; // input=3.517578125, output=-0.367189339743
			11'd901: out = 32'b10000000000000000010111101110111; // input=3.521484375, output=-0.370819912742
			11'd902: out = 32'b10000000000000000010111111101110; // input=3.525390625, output=-0.374444827485
			11'd903: out = 32'b10000000000000000011000001100100; // input=3.529296875, output=-0.378064028661
			11'd904: out = 32'b10000000000000000011000011011011; // input=3.533203125, output=-0.381677461046
			11'd905: out = 32'b10000000000000000011000101010001; // input=3.537109375, output=-0.385285069501
			11'd906: out = 32'b10000000000000000011000111000111; // input=3.541015625, output=-0.388886798981
			11'd907: out = 32'b10000000000000000011001000111101; // input=3.544921875, output=-0.392482594526
			11'd908: out = 32'b10000000000000000011001010110011; // input=3.548828125, output=-0.39607240127
			11'd909: out = 32'b10000000000000000011001100101000; // input=3.552734375, output=-0.399656164437
			11'd910: out = 32'b10000000000000000011001110011101; // input=3.556640625, output=-0.403233829342
			11'd911: out = 32'b10000000000000000011010000010010; // input=3.560546875, output=-0.406805341395
			11'd912: out = 32'b10000000000000000011010010000111; // input=3.564453125, output=-0.410370646099
			11'd913: out = 32'b10000000000000000011010011111100; // input=3.568359375, output=-0.413929689052
			11'd914: out = 32'b10000000000000000011010101110000; // input=3.572265625, output=-0.417482415947
			11'd915: out = 32'b10000000000000000011010111100100; // input=3.576171875, output=-0.421028772574
			11'd916: out = 32'b10000000000000000011011001011000; // input=3.580078125, output=-0.42456870482
			11'd917: out = 32'b10000000000000000011011011001100; // input=3.583984375, output=-0.42810215867
			11'd918: out = 32'b10000000000000000011011101000000; // input=3.587890625, output=-0.431629080208
			11'd919: out = 32'b10000000000000000011011110110011; // input=3.591796875, output=-0.435149415617
			11'd920: out = 32'b10000000000000000011100000100110; // input=3.595703125, output=-0.438663111181
			11'd921: out = 32'b10000000000000000011100010011001; // input=3.599609375, output=-0.442170113286
			11'd922: out = 32'b10000000000000000011100100001100; // input=3.603515625, output=-0.445670368419
			11'd923: out = 32'b10000000000000000011100101111110; // input=3.607421875, output=-0.44916382317
			11'd924: out = 32'b10000000000000000011100111110000; // input=3.611328125, output=-0.452650424234
			11'd925: out = 32'b10000000000000000011101001100010; // input=3.615234375, output=-0.45613011841
			11'd926: out = 32'b10000000000000000011101011010100; // input=3.619140625, output=-0.459602852601
			11'd927: out = 32'b10000000000000000011101101000110; // input=3.623046875, output=-0.463068573818
			11'd928: out = 32'b10000000000000000011101110110111; // input=3.626953125, output=-0.466527229179
			11'd929: out = 32'b10000000000000000011110000101000; // input=3.630859375, output=-0.469978765908
			11'd930: out = 32'b10000000000000000011110010011001; // input=3.634765625, output=-0.473423131339
			11'd931: out = 32'b10000000000000000011110100001010; // input=3.638671875, output=-0.476860272915
			11'd932: out = 32'b10000000000000000011110101111010; // input=3.642578125, output=-0.480290138191
			11'd933: out = 32'b10000000000000000011110111101010; // input=3.646484375, output=-0.48371267483
			11'd934: out = 32'b10000000000000000011111001011010; // input=3.650390625, output=-0.487127830609
			11'd935: out = 32'b10000000000000000011111011001010; // input=3.654296875, output=-0.490535553416
			11'd936: out = 32'b10000000000000000011111100111001; // input=3.658203125, output=-0.493935791254
			11'd937: out = 32'b10000000000000000011111110101000; // input=3.662109375, output=-0.49732849224
			11'd938: out = 32'b10000000000000000100000000010111; // input=3.666015625, output=-0.500713604605
			11'd939: out = 32'b10000000000000000100000010000110; // input=3.669921875, output=-0.504091076697
			11'd940: out = 32'b10000000000000000100000011110100; // input=3.673828125, output=-0.507460856978
			11'd941: out = 32'b10000000000000000100000101100011; // input=3.677734375, output=-0.510822894032
			11'd942: out = 32'b10000000000000000100000111010001; // input=3.681640625, output=-0.514177136557
			11'd943: out = 32'b10000000000000000100001000111110; // input=3.685546875, output=-0.517523533371
			11'd944: out = 32'b10000000000000000100001010101100; // input=3.689453125, output=-0.520862033412
			11'd945: out = 32'b10000000000000000100001100011001; // input=3.693359375, output=-0.52419258574
			11'd946: out = 32'b10000000000000000100001110000110; // input=3.697265625, output=-0.527515139534
			11'd947: out = 32'b10000000000000000100001111110010; // input=3.701171875, output=-0.530829644096
			11'd948: out = 32'b10000000000000000100010001011111; // input=3.705078125, output=-0.534136048851
			11'd949: out = 32'b10000000000000000100010011001011; // input=3.708984375, output=-0.537434303347
			11'd950: out = 32'b10000000000000000100010100110110; // input=3.712890625, output=-0.540724357256
			11'd951: out = 32'b10000000000000000100010110100010; // input=3.716796875, output=-0.544006160377
			11'd952: out = 32'b10000000000000000100011000001101; // input=3.720703125, output=-0.547279662634
			11'd953: out = 32'b10000000000000000100011001111000; // input=3.724609375, output=-0.550544814076
			11'd954: out = 32'b10000000000000000100011011100011; // input=3.728515625, output=-0.553801564881
			11'd955: out = 32'b10000000000000000100011101001101; // input=3.732421875, output=-0.557049865356
			11'd956: out = 32'b10000000000000000100011110111000; // input=3.736328125, output=-0.560289665936
			11'd957: out = 32'b10000000000000000100100000100001; // input=3.740234375, output=-0.563520917184
			11'd958: out = 32'b10000000000000000100100010001011; // input=3.744140625, output=-0.566743569797
			11'd959: out = 32'b10000000000000000100100011110100; // input=3.748046875, output=-0.5699575746
			11'd960: out = 32'b10000000000000000100100101011101; // input=3.751953125, output=-0.573162882552
			11'd961: out = 32'b10000000000000000100100111000110; // input=3.755859375, output=-0.576359444743
			11'd962: out = 32'b10000000000000000100101000101111; // input=3.759765625, output=-0.579547212398
			11'd963: out = 32'b10000000000000000100101010010111; // input=3.763671875, output=-0.582726136876
			11'd964: out = 32'b10000000000000000100101011111111; // input=3.767578125, output=-0.58589616967
			11'd965: out = 32'b10000000000000000100101101100110; // input=3.771484375, output=-0.58905726241
			11'd966: out = 32'b10000000000000000100101111001110; // input=3.775390625, output=-0.59220936686
			11'd967: out = 32'b10000000000000000100110000110101; // input=3.779296875, output=-0.595352434924
			11'd968: out = 32'b10000000000000000100110010011011; // input=3.783203125, output=-0.598486418642
			11'd969: out = 32'b10000000000000000100110100000010; // input=3.787109375, output=-0.601611270194
			11'd970: out = 32'b10000000000000000100110101101000; // input=3.791015625, output=-0.604726941898
			11'd971: out = 32'b10000000000000000100110111001101; // input=3.794921875, output=-0.607833386213
			11'd972: out = 32'b10000000000000000100111000110011; // input=3.798828125, output=-0.610930555738
			11'd973: out = 32'b10000000000000000100111010011000; // input=3.802734375, output=-0.614018403215
			11'd974: out = 32'b10000000000000000100111011111101; // input=3.806640625, output=-0.617096881526
			11'd975: out = 32'b10000000000000000100111101100010; // input=3.810546875, output=-0.620165943698
			11'd976: out = 32'b10000000000000000100111111000110; // input=3.814453125, output=-0.623225542901
			11'd977: out = 32'b10000000000000000101000000101010; // input=3.818359375, output=-0.626275632449
			11'd978: out = 32'b10000000000000000101000010001101; // input=3.822265625, output=-0.629316165801
			11'd979: out = 32'b10000000000000000101000011110001; // input=3.826171875, output=-0.632347096563
			11'd980: out = 32'b10000000000000000101000101010100; // input=3.830078125, output=-0.635368378486
			11'd981: out = 32'b10000000000000000101000110110110; // input=3.833984375, output=-0.638379965469
			11'd982: out = 32'b10000000000000000101001000011001; // input=3.837890625, output=-0.64138181156
			11'd983: out = 32'b10000000000000000101001001111011; // input=3.841796875, output=-0.644373870953
			11'd984: out = 32'b10000000000000000101001011011101; // input=3.845703125, output=-0.647356097993
			11'd985: out = 32'b10000000000000000101001100111110; // input=3.849609375, output=-0.650328447176
			11'd986: out = 32'b10000000000000000101001110011111; // input=3.853515625, output=-0.653290873148
			11'd987: out = 32'b10000000000000000101010000000000; // input=3.857421875, output=-0.656243330704
			11'd988: out = 32'b10000000000000000101010001100000; // input=3.861328125, output=-0.659185774794
			11'd989: out = 32'b10000000000000000101010011000000; // input=3.865234375, output=-0.662118160521
			11'd990: out = 32'b10000000000000000101010100100000; // input=3.869140625, output=-0.665040443139
			11'd991: out = 32'b10000000000000000101010101111111; // input=3.873046875, output=-0.667952578058
			11'd992: out = 32'b10000000000000000101010111011111; // input=3.876953125, output=-0.670854520842
			11'd993: out = 32'b10000000000000000101011000111101; // input=3.880859375, output=-0.673746227212
			11'd994: out = 32'b10000000000000000101011010011100; // input=3.884765625, output=-0.676627653043
			11'd995: out = 32'b10000000000000000101011011111010; // input=3.888671875, output=-0.679498754369
			11'd996: out = 32'b10000000000000000101011101011000; // input=3.892578125, output=-0.68235948738
			11'd997: out = 32'b10000000000000000101011110110101; // input=3.896484375, output=-0.685209808425
			11'd998: out = 32'b10000000000000000101100000010010; // input=3.900390625, output=-0.688049674011
			11'd999: out = 32'b10000000000000000101100001101111; // input=3.904296875, output=-0.690879040805
			11'd1000: out = 32'b10000000000000000101100011001011; // input=3.908203125, output=-0.693697865636
			11'd1001: out = 32'b10000000000000000101100100100111; // input=3.912109375, output=-0.69650610549
			11'd1002: out = 32'b10000000000000000101100110000011; // input=3.916015625, output=-0.699303717518
			11'd1003: out = 32'b10000000000000000101100111011110; // input=3.919921875, output=-0.702090659032
			11'd1004: out = 32'b10000000000000000101101000111001; // input=3.923828125, output=-0.704866887506
			11'd1005: out = 32'b10000000000000000101101010010100; // input=3.927734375, output=-0.707632360579
			11'd1006: out = 32'b10000000000000000101101011101110; // input=3.931640625, output=-0.710387036053
			11'd1007: out = 32'b10000000000000000101101101001000; // input=3.935546875, output=-0.713130871894
			11'd1008: out = 32'b10000000000000000101101110100001; // input=3.939453125, output=-0.715863826236
			11'd1009: out = 32'b10000000000000000101101111111011; // input=3.943359375, output=-0.718585857376
			11'd1010: out = 32'b10000000000000000101110001010011; // input=3.947265625, output=-0.72129692378
			11'd1011: out = 32'b10000000000000000101110010101100; // input=3.951171875, output=-0.723996984081
			11'd1012: out = 32'b10000000000000000101110100000100; // input=3.955078125, output=-0.726685997079
			11'd1013: out = 32'b10000000000000000101110101011100; // input=3.958984375, output=-0.729363921742
			11'd1014: out = 32'b10000000000000000101110110110011; // input=3.962890625, output=-0.732030717209
			11'd1015: out = 32'b10000000000000000101111000001010; // input=3.966796875, output=-0.734686342788
			11'd1016: out = 32'b10000000000000000101111001100001; // input=3.970703125, output=-0.737330757958
			11'd1017: out = 32'b10000000000000000101111010110111; // input=3.974609375, output=-0.739963922367
			11'd1018: out = 32'b10000000000000000101111100001101; // input=3.978515625, output=-0.742585795837
			11'd1019: out = 32'b10000000000000000101111101100011; // input=3.982421875, output=-0.745196338362
			11'd1020: out = 32'b10000000000000000101111110111000; // input=3.986328125, output=-0.747795510107
			11'd1021: out = 32'b10000000000000000110000000001101; // input=3.990234375, output=-0.750383271413
			11'd1022: out = 32'b10000000000000000110000001100001; // input=3.994140625, output=-0.752959582793
			11'd1023: out = 32'b10000000000000000110000010110101; // input=3.998046875, output=-0.755524404937
			11'd1024: out = 32'b10000000000000000000000001000000; // input=-0.001953125, output=-0.00195312375824
			11'd1025: out = 32'b10000000000000000000000011000000; // input=-0.005859375, output=-0.00585934147244
			11'd1026: out = 32'b10000000000000000000000101000000; // input=-0.009765625, output=-0.00976546978031
			11'd1027: out = 32'b10000000000000000000000111000000; // input=-0.013671875, output=-0.0136714490791
			11'd1028: out = 32'b10000000000000000000001001000000; // input=-0.017578125, output=-0.0175772197684
			11'd1029: out = 32'b10000000000000000000001011000000; // input=-0.021484375, output=-0.021482722251
			11'd1030: out = 32'b10000000000000000000001101000000; // input=-0.025390625, output=-0.0253878969337
			11'd1031: out = 32'b10000000000000000000001111000000; // input=-0.029296875, output=-0.0292926842283
			11'd1032: out = 32'b10000000000000000000010001000000; // input=-0.033203125, output=-0.0331970245525
			11'd1033: out = 32'b10000000000000000000010011000000; // input=-0.037109375, output=-0.0371008583311
			11'd1034: out = 32'b10000000000000000000010101000000; // input=-0.041015625, output=-0.0410041259961
			11'd1035: out = 32'b10000000000000000000010111000000; // input=-0.044921875, output=-0.0449067679887
			11'd1036: out = 32'b10000000000000000000011000111111; // input=-0.048828125, output=-0.0488087247592
			11'd1037: out = 32'b10000000000000000000011010111111; // input=-0.052734375, output=-0.0527099367686
			11'd1038: out = 32'b10000000000000000000011100111111; // input=-0.056640625, output=-0.0566103444893
			11'd1039: out = 32'b10000000000000000000011110111111; // input=-0.060546875, output=-0.0605098884057
			11'd1040: out = 32'b10000000000000000000100000111111; // input=-0.064453125, output=-0.0644085090157
			11'd1041: out = 32'b10000000000000000000100010111110; // input=-0.068359375, output=-0.0683061468311
			11'd1042: out = 32'b10000000000000000000100100111110; // input=-0.072265625, output=-0.0722027423787
			11'd1043: out = 32'b10000000000000000000100110111110; // input=-0.076171875, output=-0.0760982362014
			11'd1044: out = 32'b10000000000000000000101000111101; // input=-0.080078125, output=-0.0799925688585
			11'd1045: out = 32'b10000000000000000000101010111101; // input=-0.083984375, output=-0.0838856809275
			11'd1046: out = 32'b10000000000000000000101100111100; // input=-0.087890625, output=-0.0877775130042
			11'd1047: out = 32'b10000000000000000000101110111100; // input=-0.091796875, output=-0.091668005704
			11'd1048: out = 32'b10000000000000000000110000111011; // input=-0.095703125, output=-0.0955570996629
			11'd1049: out = 32'b10000000000000000000110010111011; // input=-0.099609375, output=-0.099444735538
			11'd1050: out = 32'b10000000000000000000110100111010; // input=-0.103515625, output=-0.103330854009
			11'd1051: out = 32'b10000000000000000000110110111001; // input=-0.107421875, output=-0.107215395778
			11'd1052: out = 32'b10000000000000000000111000111000; // input=-0.111328125, output=-0.111098301572
			11'd1053: out = 32'b10000000000000000000111010111000; // input=-0.115234375, output=-0.114979512142
			11'd1054: out = 32'b10000000000000000000111100110111; // input=-0.119140625, output=-0.118858968267
			11'd1055: out = 32'b10000000000000000000111110110110; // input=-0.123046875, output=-0.12273661075
			11'd1056: out = 32'b10000000000000000001000000110101; // input=-0.126953125, output=-0.126612380424
			11'd1057: out = 32'b10000000000000000001000010110100; // input=-0.130859375, output=-0.130486218148
			11'd1058: out = 32'b10000000000000000001000100110011; // input=-0.134765625, output=-0.134358064813
			11'd1059: out = 32'b10000000000000000001000110110001; // input=-0.138671875, output=-0.13822786134
			11'd1060: out = 32'b10000000000000000001001000110000; // input=-0.142578125, output=-0.142095548679
			11'd1061: out = 32'b10000000000000000001001010101111; // input=-0.146484375, output=-0.145961067815
			11'd1062: out = 32'b10000000000000000001001100101101; // input=-0.150390625, output=-0.149824359765
			11'd1063: out = 32'b10000000000000000001001110101100; // input=-0.154296875, output=-0.153685365579
			11'd1064: out = 32'b10000000000000000001010000101010; // input=-0.158203125, output=-0.157544026344
			11'd1065: out = 32'b10000000000000000001010010101001; // input=-0.162109375, output=-0.161400283181
			11'd1066: out = 32'b10000000000000000001010100100111; // input=-0.166015625, output=-0.165254077248
			11'd1067: out = 32'b10000000000000000001010110100101; // input=-0.169921875, output=-0.169105349741
			11'd1068: out = 32'b10000000000000000001011000100011; // input=-0.173828125, output=-0.172954041894
			11'd1069: out = 32'b10000000000000000001011010100001; // input=-0.177734375, output=-0.176800094982
			11'd1070: out = 32'b10000000000000000001011100011111; // input=-0.181640625, output=-0.180643450318
			11'd1071: out = 32'b10000000000000000001011110011101; // input=-0.185546875, output=-0.184484049257
			11'd1072: out = 32'b10000000000000000001100000011011; // input=-0.189453125, output=-0.188321833196
			11'd1073: out = 32'b10000000000000000001100010011001; // input=-0.193359375, output=-0.192156743576
			11'd1074: out = 32'b10000000000000000001100100010110; // input=-0.197265625, output=-0.19598872188
			11'd1075: out = 32'b10000000000000000001100110010100; // input=-0.201171875, output=-0.199817709638
			11'd1076: out = 32'b10000000000000000001101000010001; // input=-0.205078125, output=-0.203643648423
			11'd1077: out = 32'b10000000000000000001101010001110; // input=-0.208984375, output=-0.207466479857
			11'd1078: out = 32'b10000000000000000001101100001011; // input=-0.212890625, output=-0.211286145607
			11'd1079: out = 32'b10000000000000000001101110001000; // input=-0.216796875, output=-0.215102587391
			11'd1080: out = 32'b10000000000000000001110000000101; // input=-0.220703125, output=-0.218915746974
			11'd1081: out = 32'b10000000000000000001110010000010; // input=-0.224609375, output=-0.222725566172
			11'd1082: out = 32'b10000000000000000001110011111111; // input=-0.228515625, output=-0.226531986852
			11'd1083: out = 32'b10000000000000000001110101111100; // input=-0.232421875, output=-0.230334950932
			11'd1084: out = 32'b10000000000000000001110111111000; // input=-0.236328125, output=-0.234134400385
			11'd1085: out = 32'b10000000000000000001111001110100; // input=-0.240234375, output=-0.237930277234
			11'd1086: out = 32'b10000000000000000001111011110001; // input=-0.244140625, output=-0.241722523561
			11'd1087: out = 32'b10000000000000000001111101101101; // input=-0.248046875, output=-0.245511081499
			11'd1088: out = 32'b10000000000000000001111111101001; // input=-0.251953125, output=-0.24929589324
			11'd1089: out = 32'b10000000000000000010000001100101; // input=-0.255859375, output=-0.253076901032
			11'd1090: out = 32'b10000000000000000010000011100001; // input=-0.259765625, output=-0.256854047182
			11'd1091: out = 32'b10000000000000000010000101011100; // input=-0.263671875, output=-0.260627274056
			11'd1092: out = 32'b10000000000000000010000111011000; // input=-0.267578125, output=-0.264396524078
			11'd1093: out = 32'b10000000000000000010001001010011; // input=-0.271484375, output=-0.268161739734
			11'd1094: out = 32'b10000000000000000010001011001110; // input=-0.275390625, output=-0.271922863572
			11'd1095: out = 32'b10000000000000000010001101001001; // input=-0.279296875, output=-0.275679838202
			11'd1096: out = 32'b10000000000000000010001111000100; // input=-0.283203125, output=-0.279432606296
			11'd1097: out = 32'b10000000000000000010010000111111; // input=-0.287109375, output=-0.283181110593
			11'd1098: out = 32'b10000000000000000010010010111010; // input=-0.291015625, output=-0.286925293895
			11'd1099: out = 32'b10000000000000000010010100110101; // input=-0.294921875, output=-0.290665099069
			11'd1100: out = 32'b10000000000000000010010110101111; // input=-0.298828125, output=-0.294400469052
			11'd1101: out = 32'b10000000000000000010011000101001; // input=-0.302734375, output=-0.298131346846
			11'd1102: out = 32'b10000000000000000010011010100011; // input=-0.306640625, output=-0.301857675522
			11'd1103: out = 32'b10000000000000000010011100011101; // input=-0.310546875, output=-0.305579398221
			11'd1104: out = 32'b10000000000000000010011110010111; // input=-0.314453125, output=-0.309296458155
			11'd1105: out = 32'b10000000000000000010100000010001; // input=-0.318359375, output=-0.313008798605
			11'd1106: out = 32'b10000000000000000010100010001010; // input=-0.322265625, output=-0.316716362927
			11'd1107: out = 32'b10000000000000000010100100000011; // input=-0.326171875, output=-0.320419094546
			11'd1108: out = 32'b10000000000000000010100101111101; // input=-0.330078125, output=-0.324116936964
			11'd1109: out = 32'b10000000000000000010100111110110; // input=-0.333984375, output=-0.327809833756
			11'd1110: out = 32'b10000000000000000010101001101111; // input=-0.337890625, output=-0.331497728574
			11'd1111: out = 32'b10000000000000000010101011100111; // input=-0.341796875, output=-0.335180565144
			11'd1112: out = 32'b10000000000000000010101101100000; // input=-0.345703125, output=-0.338858287271
			11'd1113: out = 32'b10000000000000000010101111011000; // input=-0.349609375, output=-0.342530838838
			11'd1114: out = 32'b10000000000000000010110001010000; // input=-0.353515625, output=-0.346198163805
			11'd1115: out = 32'b10000000000000000010110011001000; // input=-0.357421875, output=-0.349860206215
			11'd1116: out = 32'b10000000000000000010110101000000; // input=-0.361328125, output=-0.353516910188
			11'd1117: out = 32'b10000000000000000010110110111000; // input=-0.365234375, output=-0.357168219928
			11'd1118: out = 32'b10000000000000000010111000101111; // input=-0.369140625, output=-0.36081407972
			11'd1119: out = 32'b10000000000000000010111010100110; // input=-0.373046875, output=-0.364454433933
			11'd1120: out = 32'b10000000000000000010111100011110; // input=-0.376953125, output=-0.36808922702
			11'd1121: out = 32'b10000000000000000010111110010100; // input=-0.380859375, output=-0.371718403519
			11'd1122: out = 32'b10000000000000000011000000001011; // input=-0.384765625, output=-0.375341908052
			11'd1123: out = 32'b10000000000000000011000010000010; // input=-0.388671875, output=-0.378959685329
			11'd1124: out = 32'b10000000000000000011000011111000; // input=-0.392578125, output=-0.382571680148
			11'd1125: out = 32'b10000000000000000011000101101110; // input=-0.396484375, output=-0.386177837393
			11'd1126: out = 32'b10000000000000000011000111100100; // input=-0.400390625, output=-0.38977810204
			11'd1127: out = 32'b10000000000000000011001001011010; // input=-0.404296875, output=-0.393372419153
			11'd1128: out = 32'b10000000000000000011001011010000; // input=-0.408203125, output=-0.396960733886
			11'd1129: out = 32'b10000000000000000011001101000101; // input=-0.412109375, output=-0.400542991487
			11'd1130: out = 32'b10000000000000000011001110111010; // input=-0.416015625, output=-0.404119137295
			11'd1131: out = 32'b10000000000000000011010000101111; // input=-0.419921875, output=-0.407689116742
			11'd1132: out = 32'b10000000000000000011010010100100; // input=-0.423828125, output=-0.411252875354
			11'd1133: out = 32'b10000000000000000011010100011001; // input=-0.427734375, output=-0.414810358754
			11'd1134: out = 32'b10000000000000000011010110001101; // input=-0.431640625, output=-0.418361512658
			11'd1135: out = 32'b10000000000000000011011000000001; // input=-0.435546875, output=-0.42190628288
			11'd1136: out = 32'b10000000000000000011011001110101; // input=-0.439453125, output=-0.425444615332
			11'd1137: out = 32'b10000000000000000011011011101001; // input=-0.443359375, output=-0.428976456021
			11'd1138: out = 32'b10000000000000000011011101011100; // input=-0.447265625, output=-0.432501751058
			11'd1139: out = 32'b10000000000000000011011111010000; // input=-0.451171875, output=-0.436020446651
			11'd1140: out = 32'b10000000000000000011100001000011; // input=-0.455078125, output=-0.439532489107
			11'd1141: out = 32'b10000000000000000011100010110101; // input=-0.458984375, output=-0.443037824839
			11'd1142: out = 32'b10000000000000000011100100101000; // input=-0.462890625, output=-0.446536400359
			11'd1143: out = 32'b10000000000000000011100110011011; // input=-0.466796875, output=-0.450028162283
			11'd1144: out = 32'b10000000000000000011101000001101; // input=-0.470703125, output=-0.45351305733
			11'd1145: out = 32'b10000000000000000011101001111111; // input=-0.474609375, output=-0.456991032326
			11'd1146: out = 32'b10000000000000000011101011110000; // input=-0.478515625, output=-0.460462034202
			11'd1147: out = 32'b10000000000000000011101101100010; // input=-0.482421875, output=-0.463926009993
			11'd1148: out = 32'b10000000000000000011101111010011; // input=-0.486328125, output=-0.467382906844
			11'd1149: out = 32'b10000000000000000011110001000100; // input=-0.490234375, output=-0.470832672007
			11'd1150: out = 32'b10000000000000000011110010110101; // input=-0.494140625, output=-0.474275252843
			11'd1151: out = 32'b10000000000000000011110100100110; // input=-0.498046875, output=-0.477710596821
			11'd1152: out = 32'b10000000000000000011110110010110; // input=-0.501953125, output=-0.481138651524
			11'd1153: out = 32'b10000000000000000011111000000110; // input=-0.505859375, output=-0.484559364643
			11'd1154: out = 32'b10000000000000000011111001110110; // input=-0.509765625, output=-0.487972683983
			11'd1155: out = 32'b10000000000000000011111011100101; // input=-0.513671875, output=-0.491378557459
			11'd1156: out = 32'b10000000000000000011111101010101; // input=-0.517578125, output=-0.494776933103
			11'd1157: out = 32'b10000000000000000011111111000100; // input=-0.521484375, output=-0.49816775906
			11'd1158: out = 32'b10000000000000000100000000110011; // input=-0.525390625, output=-0.50155098359
			11'd1159: out = 32'b10000000000000000100000010100001; // input=-0.529296875, output=-0.504926555069
			11'd1160: out = 32'b10000000000000000100000100010000; // input=-0.533203125, output=-0.50829442199
			11'd1161: out = 32'b10000000000000000100000101111110; // input=-0.537109375, output=-0.511654532964
			11'd1162: out = 32'b10000000000000000100000111101100; // input=-0.541015625, output=-0.515006836719
			11'd1163: out = 32'b10000000000000000100001001011001; // input=-0.544921875, output=-0.518351282103
			11'd1164: out = 32'b10000000000000000100001011000111; // input=-0.548828125, output=-0.521687818084
			11'd1165: out = 32'b10000000000000000100001100110100; // input=-0.552734375, output=-0.525016393751
			11'd1166: out = 32'b10000000000000000100001110100001; // input=-0.556640625, output=-0.528336958314
			11'd1167: out = 32'b10000000000000000100010000001101; // input=-0.560546875, output=-0.531649461105
			11'd1168: out = 32'b10000000000000000100010001111001; // input=-0.564453125, output=-0.534953851579
			11'd1169: out = 32'b10000000000000000100010011100101; // input=-0.568359375, output=-0.538250079316
			11'd1170: out = 32'b10000000000000000100010101010001; // input=-0.572265625, output=-0.541538094019
			11'd1171: out = 32'b10000000000000000100010110111101; // input=-0.576171875, output=-0.544817845516
			11'd1172: out = 32'b10000000000000000100011000101000; // input=-0.580078125, output=-0.548089283764
			11'd1173: out = 32'b10000000000000000100011010010011; // input=-0.583984375, output=-0.551352358843
			11'd1174: out = 32'b10000000000000000100011011111101; // input=-0.587890625, output=-0.554607020964
			11'd1175: out = 32'b10000000000000000100011101101000; // input=-0.591796875, output=-0.557853220464
			11'd1176: out = 32'b10000000000000000100011111010010; // input=-0.595703125, output=-0.561090907811
			11'd1177: out = 32'b10000000000000000100100000111100; // input=-0.599609375, output=-0.5643200336
			11'd1178: out = 32'b10000000000000000100100010100101; // input=-0.603515625, output=-0.56754054856
			11'd1179: out = 32'b10000000000000000100100100001110; // input=-0.607421875, output=-0.570752403549
			11'd1180: out = 32'b10000000000000000100100101110111; // input=-0.611328125, output=-0.573955549559
			11'd1181: out = 32'b10000000000000000100100111100000; // input=-0.615234375, output=-0.577149937714
			11'd1182: out = 32'b10000000000000000100101001001000; // input=-0.619140625, output=-0.58033551927
			11'd1183: out = 32'b10000000000000000100101010110001; // input=-0.623046875, output=-0.583512245621
			11'd1184: out = 32'b10000000000000000100101100011000; // input=-0.626953125, output=-0.586680068292
			11'd1185: out = 32'b10000000000000000100101110000000; // input=-0.630859375, output=-0.589838938948
			11'd1186: out = 32'b10000000000000000100101111100111; // input=-0.634765625, output=-0.592988809387
			11'd1187: out = 32'b10000000000000000100110001001110; // input=-0.638671875, output=-0.596129631546
			11'd1188: out = 32'b10000000000000000100110010110101; // input=-0.642578125, output=-0.599261357501
			11'd1189: out = 32'b10000000000000000100110100011011; // input=-0.646484375, output=-0.602383939464
			11'd1190: out = 32'b10000000000000000100110110000001; // input=-0.650390625, output=-0.60549732979
			11'd1191: out = 32'b10000000000000000100110111100111; // input=-0.654296875, output=-0.608601480971
			11'd1192: out = 32'b10000000000000000100111001001100; // input=-0.658203125, output=-0.611696345643
			11'd1193: out = 32'b10000000000000000100111010110001; // input=-0.662109375, output=-0.614781876581
			11'd1194: out = 32'b10000000000000000100111100010110; // input=-0.666015625, output=-0.617858026704
			11'd1195: out = 32'b10000000000000000100111101111010; // input=-0.669921875, output=-0.620924749074
			11'd1196: out = 32'b10000000000000000100111111011111; // input=-0.673828125, output=-0.623981996896
			11'd1197: out = 32'b10000000000000000101000001000011; // input=-0.677734375, output=-0.62702972352
			11'd1198: out = 32'b10000000000000000101000010100110; // input=-0.681640625, output=-0.630067882443
			11'd1199: out = 32'b10000000000000000101000100001001; // input=-0.685546875, output=-0.633096427304
			11'd1200: out = 32'b10000000000000000101000101101100; // input=-0.689453125, output=-0.636115311893
			11'd1201: out = 32'b10000000000000000101000111001111; // input=-0.693359375, output=-0.639124490145
			11'd1202: out = 32'b10000000000000000101001000110001; // input=-0.697265625, output=-0.642123916144
			11'd1203: out = 32'b10000000000000000101001010010011; // input=-0.701171875, output=-0.645113544122
			11'd1204: out = 32'b10000000000000000101001011110101; // input=-0.705078125, output=-0.64809332846
			11'd1205: out = 32'b10000000000000000101001101010110; // input=-0.708984375, output=-0.651063223692
			11'd1206: out = 32'b10000000000000000101001110110111; // input=-0.712890625, output=-0.6540231845
			11'd1207: out = 32'b10000000000000000101010000011000; // input=-0.716796875, output=-0.65697316572
			11'd1208: out = 32'b10000000000000000101010001111000; // input=-0.720703125, output=-0.659913122336
			11'd1209: out = 32'b10000000000000000101010011011000; // input=-0.724609375, output=-0.662843009491
			11'd1210: out = 32'b10000000000000000101010100111000; // input=-0.728515625, output=-0.665762782477
			11'd1211: out = 32'b10000000000000000101010110010111; // input=-0.732421875, output=-0.668672396741
			11'd1212: out = 32'b10000000000000000101010111110110; // input=-0.736328125, output=-0.671571807888
			11'd1213: out = 32'b10000000000000000101011001010101; // input=-0.740234375, output=-0.674460971675
			11'd1214: out = 32'b10000000000000000101011010110011; // input=-0.744140625, output=-0.677339844018
			11'd1215: out = 32'b10000000000000000101011100010001; // input=-0.748046875, output=-0.680208380988
			11'd1216: out = 32'b10000000000000000101011101101111; // input=-0.751953125, output=-0.683066538814
			11'd1217: out = 32'b10000000000000000101011111001100; // input=-0.755859375, output=-0.685914273886
			11'd1218: out = 32'b10000000000000000101100000101001; // input=-0.759765625, output=-0.68875154275
			11'd1219: out = 32'b10000000000000000101100010000110; // input=-0.763671875, output=-0.691578302113
			11'd1220: out = 32'b10000000000000000101100011100010; // input=-0.767578125, output=-0.694394508842
			11'd1221: out = 32'b10000000000000000101100100111110; // input=-0.771484375, output=-0.697200119965
			11'd1222: out = 32'b10000000000000000101100110011001; // input=-0.775390625, output=-0.699995092672
			11'd1223: out = 32'b10000000000000000101100111110101; // input=-0.779296875, output=-0.702779384315
			11'd1224: out = 32'b10000000000000000101101001010000; // input=-0.783203125, output=-0.705552952409
			11'd1225: out = 32'b10000000000000000101101010101010; // input=-0.787109375, output=-0.708315754633
			11'd1226: out = 32'b10000000000000000101101100000100; // input=-0.791015625, output=-0.711067748831
			11'd1227: out = 32'b10000000000000000101101101011110; // input=-0.794921875, output=-0.713808893009
			11'd1228: out = 32'b10000000000000000101101110111000; // input=-0.798828125, output=-0.716539145342
			11'd1229: out = 32'b10000000000000000101110000010001; // input=-0.802734375, output=-0.719258464169
			11'd1230: out = 32'b10000000000000000101110001101001; // input=-0.806640625, output=-0.721966807997
			11'd1231: out = 32'b10000000000000000101110011000010; // input=-0.810546875, output=-0.7246641355
			11'd1232: out = 32'b10000000000000000101110100011010; // input=-0.814453125, output=-0.727350405519
			11'd1233: out = 32'b10000000000000000101110101110001; // input=-0.818359375, output=-0.730025577067
			11'd1234: out = 32'b10000000000000000101110111001001; // input=-0.822265625, output=-0.732689609322
			11'd1235: out = 32'b10000000000000000101111000100000; // input=-0.826171875, output=-0.735342461635
			11'd1236: out = 32'b10000000000000000101111001110110; // input=-0.830078125, output=-0.737984093527
			11'd1237: out = 32'b10000000000000000101111011001100; // input=-0.833984375, output=-0.740614464689
			11'd1238: out = 32'b10000000000000000101111100100010; // input=-0.837890625, output=-0.743233534986
			11'd1239: out = 32'b10000000000000000101111101111000; // input=-0.841796875, output=-0.745841264454
			11'd1240: out = 32'b10000000000000000101111111001101; // input=-0.845703125, output=-0.748437613302
			11'd1241: out = 32'b10000000000000000110000000100010; // input=-0.849609375, output=-0.751022541912
			11'd1242: out = 32'b10000000000000000110000001110110; // input=-0.853515625, output=-0.753596010843
			11'd1243: out = 32'b10000000000000000110000011001010; // input=-0.857421875, output=-0.756157980826
			11'd1244: out = 32'b10000000000000000110000100011101; // input=-0.861328125, output=-0.758708412768
			11'd1245: out = 32'b10000000000000000110000101110001; // input=-0.865234375, output=-0.761247267753
			11'd1246: out = 32'b10000000000000000110000111000011; // input=-0.869140625, output=-0.763774507042
			11'd1247: out = 32'b10000000000000000110001000010110; // input=-0.873046875, output=-0.766290092071
			11'd1248: out = 32'b10000000000000000110001001101000; // input=-0.876953125, output=-0.768793984456
			11'd1249: out = 32'b10000000000000000110001010111010; // input=-0.880859375, output=-0.771286145991
			11'd1250: out = 32'b10000000000000000110001100001011; // input=-0.884765625, output=-0.773766538648
			11'd1251: out = 32'b10000000000000000110001101011100; // input=-0.888671875, output=-0.77623512458
			11'd1252: out = 32'b10000000000000000110001110101100; // input=-0.892578125, output=-0.778691866119
			11'd1253: out = 32'b10000000000000000110001111111100; // input=-0.896484375, output=-0.781136725778
			11'd1254: out = 32'b10000000000000000110010001001100; // input=-0.900390625, output=-0.783569666252
			11'd1255: out = 32'b10000000000000000110010010011011; // input=-0.904296875, output=-0.785990650417
			11'd1256: out = 32'b10000000000000000110010011101010; // input=-0.908203125, output=-0.788399641331
			11'd1257: out = 32'b10000000000000000110010100111001; // input=-0.912109375, output=-0.790796602237
			11'd1258: out = 32'b10000000000000000110010110000111; // input=-0.916015625, output=-0.79318149656
			11'd1259: out = 32'b10000000000000000110010111010101; // input=-0.919921875, output=-0.795554287909
			11'd1260: out = 32'b10000000000000000110011000100010; // input=-0.923828125, output=-0.797914940078
			11'd1261: out = 32'b10000000000000000110011001101111; // input=-0.927734375, output=-0.800263417047
			11'd1262: out = 32'b10000000000000000110011010111100; // input=-0.931640625, output=-0.802599682981
			11'd1263: out = 32'b10000000000000000110011100001000; // input=-0.935546875, output=-0.804923702231
			11'd1264: out = 32'b10000000000000000110011101010011; // input=-0.939453125, output=-0.807235439336
			11'd1265: out = 32'b10000000000000000110011110011111; // input=-0.943359375, output=-0.809534859021
			11'd1266: out = 32'b10000000000000000110011111101010; // input=-0.947265625, output=-0.8118219262
			11'd1267: out = 32'b10000000000000000110100000110100; // input=-0.951171875, output=-0.814096605976
			11'd1268: out = 32'b10000000000000000110100001111110; // input=-0.955078125, output=-0.816358863639
			11'd1269: out = 32'b10000000000000000110100011001000; // input=-0.958984375, output=-0.81860866467
			11'd1270: out = 32'b10000000000000000110100100010001; // input=-0.962890625, output=-0.82084597474
			11'd1271: out = 32'b10000000000000000110100101011010; // input=-0.966796875, output=-0.82307075971
			11'd1272: out = 32'b10000000000000000110100110100011; // input=-0.970703125, output=-0.825282985633
			11'd1273: out = 32'b10000000000000000110100111101011; // input=-0.974609375, output=-0.827482618753
			11'd1274: out = 32'b10000000000000000110101000110011; // input=-0.978515625, output=-0.829669625507
			11'd1275: out = 32'b10000000000000000110101001111010; // input=-0.982421875, output=-0.831843972523
			11'd1276: out = 32'b10000000000000000110101011000001; // input=-0.986328125, output=-0.834005626623
			11'd1277: out = 32'b10000000000000000110101100000111; // input=-0.990234375, output=-0.836154554823
			11'd1278: out = 32'b10000000000000000110101101001101; // input=-0.994140625, output=-0.838290724334
			11'd1279: out = 32'b10000000000000000110101110010011; // input=-0.998046875, output=-0.84041410256
			11'd1280: out = 32'b10000000000000000110101111011000; // input=-1.001953125, output=-0.8425246571
			11'd1281: out = 32'b10000000000000000110110000011101; // input=-1.005859375, output=-0.844622355751
			11'd1282: out = 32'b10000000000000000110110001100001; // input=-1.009765625, output=-0.846707166504
			11'd1283: out = 32'b10000000000000000110110010100101; // input=-1.013671875, output=-0.848779057547
			11'd1284: out = 32'b10000000000000000110110011101000; // input=-1.017578125, output=-0.850837997266
			11'd1285: out = 32'b10000000000000000110110100101011; // input=-1.021484375, output=-0.852883954244
			11'd1286: out = 32'b10000000000000000110110101101110; // input=-1.025390625, output=-0.854916897262
			11'd1287: out = 32'b10000000000000000110110110110000; // input=-1.029296875, output=-0.8569367953
			11'd1288: out = 32'b10000000000000000110110111110010; // input=-1.033203125, output=-0.858943617537
			11'd1289: out = 32'b10000000000000000110111000110011; // input=-1.037109375, output=-0.860937333352
			11'd1290: out = 32'b10000000000000000110111001110100; // input=-1.041015625, output=-0.862917912321
			11'd1291: out = 32'b10000000000000000110111010110101; // input=-1.044921875, output=-0.864885324225
			11'd1292: out = 32'b10000000000000000110111011110101; // input=-1.048828125, output=-0.866839539044
			11'd1293: out = 32'b10000000000000000110111100110100; // input=-1.052734375, output=-0.868780526957
			11'd1294: out = 32'b10000000000000000110111101110011; // input=-1.056640625, output=-0.870708258348
			11'd1295: out = 32'b10000000000000000110111110110010; // input=-1.060546875, output=-0.872622703803
			11'd1296: out = 32'b10000000000000000110111111110000; // input=-1.064453125, output=-0.874523834109
			11'd1297: out = 32'b10000000000000000111000000101110; // input=-1.068359375, output=-0.876411620257
			11'd1298: out = 32'b10000000000000000111000001101100; // input=-1.072265625, output=-0.878286033441
			11'd1299: out = 32'b10000000000000000111000010101001; // input=-1.076171875, output=-0.880147045062
			11'd1300: out = 32'b10000000000000000111000011100101; // input=-1.080078125, output=-0.881994626722
			11'd1301: out = 32'b10000000000000000111000100100001; // input=-1.083984375, output=-0.883828750229
			11'd1302: out = 32'b10000000000000000111000101011101; // input=-1.087890625, output=-0.885649387596
			11'd1303: out = 32'b10000000000000000111000110011000; // input=-1.091796875, output=-0.887456511044
			11'd1304: out = 32'b10000000000000000111000111010011; // input=-1.095703125, output=-0.889250092997
			11'd1305: out = 32'b10000000000000000111001000001101; // input=-1.099609375, output=-0.891030106087
			11'd1306: out = 32'b10000000000000000111001001000111; // input=-1.103515625, output=-0.892796523155
			11'd1307: out = 32'b10000000000000000111001010000001; // input=-1.107421875, output=-0.894549317246
			11'd1308: out = 32'b10000000000000000111001010111010; // input=-1.111328125, output=-0.896288461615
			11'd1309: out = 32'b10000000000000000111001011110010; // input=-1.115234375, output=-0.898013929725
			11'd1310: out = 32'b10000000000000000111001100101010; // input=-1.119140625, output=-0.899725695247
			11'd1311: out = 32'b10000000000000000111001101100010; // input=-1.123046875, output=-0.901423732062
			11'd1312: out = 32'b10000000000000000111001110011001; // input=-1.126953125, output=-0.90310801426
			11'd1313: out = 32'b10000000000000000111001111010000; // input=-1.130859375, output=-0.90477851614
			11'd1314: out = 32'b10000000000000000111010000000110; // input=-1.134765625, output=-0.906435212214
			11'd1315: out = 32'b10000000000000000111010000111100; // input=-1.138671875, output=-0.908078077202
			11'd1316: out = 32'b10000000000000000111010001110001; // input=-1.142578125, output=-0.909707086035
			11'd1317: out = 32'b10000000000000000111010010100110; // input=-1.146484375, output=-0.911322213858
			11'd1318: out = 32'b10000000000000000111010011011011; // input=-1.150390625, output=-0.912923436025
			11'd1319: out = 32'b10000000000000000111010100001111; // input=-1.154296875, output=-0.914510728103
			11'd1320: out = 32'b10000000000000000111010101000010; // input=-1.158203125, output=-0.916084065873
			11'd1321: out = 32'b10000000000000000111010101110101; // input=-1.162109375, output=-0.917643425327
			11'd1322: out = 32'b10000000000000000111010110101000; // input=-1.166015625, output=-0.919188782671
			11'd1323: out = 32'b10000000000000000111010111011010; // input=-1.169921875, output=-0.920720114326
			11'd1324: out = 32'b10000000000000000111011000001100; // input=-1.173828125, output=-0.922237396924
			11'd1325: out = 32'b10000000000000000111011000111101; // input=-1.177734375, output=-0.923740607315
			11'd1326: out = 32'b10000000000000000111011001101110; // input=-1.181640625, output=-0.92522972256
			11'd1327: out = 32'b10000000000000000111011010011110; // input=-1.185546875, output=-0.926704719938
			11'd1328: out = 32'b10000000000000000111011011001110; // input=-1.189453125, output=-0.928165576942
			11'd1329: out = 32'b10000000000000000111011011111110; // input=-1.193359375, output=-0.929612271281
			11'd1330: out = 32'b10000000000000000111011100101100; // input=-1.197265625, output=-0.931044780881
			11'd1331: out = 32'b10000000000000000111011101011011; // input=-1.201171875, output=-0.932463083883
			11'd1332: out = 32'b10000000000000000111011110001001; // input=-1.205078125, output=-0.933867158646
			11'd1333: out = 32'b10000000000000000111011110110111; // input=-1.208984375, output=-0.935256983744
			11'd1334: out = 32'b10000000000000000111011111100100; // input=-1.212890625, output=-0.936632537972
			11'd1335: out = 32'b10000000000000000111100000010000; // input=-1.216796875, output=-0.93799380034
			11'd1336: out = 32'b10000000000000000111100000111100; // input=-1.220703125, output=-0.939340750076
			11'd1337: out = 32'b10000000000000000111100001101000; // input=-1.224609375, output=-0.940673366629
			11'd1338: out = 32'b10000000000000000111100010010011; // input=-1.228515625, output=-0.941991629663
			11'd1339: out = 32'b10000000000000000111100010111110; // input=-1.232421875, output=-0.943295519063
			11'd1340: out = 32'b10000000000000000111100011101000; // input=-1.236328125, output=-0.944585014935
			11'd1341: out = 32'b10000000000000000111100100010010; // input=-1.240234375, output=-0.945860097601
			11'd1342: out = 32'b10000000000000000111100100111011; // input=-1.244140625, output=-0.947120747606
			11'd1343: out = 32'b10000000000000000111100101100100; // input=-1.248046875, output=-0.948366945714
			11'd1344: out = 32'b10000000000000000111100110001100; // input=-1.251953125, output=-0.949598672909
			11'd1345: out = 32'b10000000000000000111100110110100; // input=-1.255859375, output=-0.950815910397
			11'd1346: out = 32'b10000000000000000111100111011100; // input=-1.259765625, output=-0.952018639603
			11'd1347: out = 32'b10000000000000000111101000000011; // input=-1.263671875, output=-0.953206842177
			11'd1348: out = 32'b10000000000000000111101000101001; // input=-1.267578125, output=-0.954380499987
			11'd1349: out = 32'b10000000000000000111101001001111; // input=-1.271484375, output=-0.955539595124
			11'd1350: out = 32'b10000000000000000111101001110101; // input=-1.275390625, output=-0.956684109903
			11'd1351: out = 32'b10000000000000000111101010011010; // input=-1.279296875, output=-0.95781402686
			11'd1352: out = 32'b10000000000000000111101010111110; // input=-1.283203125, output=-0.958929328753
			11'd1353: out = 32'b10000000000000000111101011100010; // input=-1.287109375, output=-0.960029998564
			11'd1354: out = 32'b10000000000000000111101100000110; // input=-1.291015625, output=-0.961116019499
			11'd1355: out = 32'b10000000000000000111101100101001; // input=-1.294921875, output=-0.962187374985
			11'd1356: out = 32'b10000000000000000111101101001100; // input=-1.298828125, output=-0.963244048676
			11'd1357: out = 32'b10000000000000000111101101101110; // input=-1.302734375, output=-0.964286024448
			11'd1358: out = 32'b10000000000000000111101110001111; // input=-1.306640625, output=-0.965313286402
			11'd1359: out = 32'b10000000000000000111101110110001; // input=-1.310546875, output=-0.966325818863
			11'd1360: out = 32'b10000000000000000111101111010001; // input=-1.314453125, output=-0.96732360638
			11'd1361: out = 32'b10000000000000000111101111110001; // input=-1.318359375, output=-0.96830663373
			11'd1362: out = 32'b10000000000000000111110000010001; // input=-1.322265625, output=-0.969274885911
			11'd1363: out = 32'b10000000000000000111110000110000; // input=-1.326171875, output=-0.970228348151
			11'd1364: out = 32'b10000000000000000111110001001111; // input=-1.330078125, output=-0.971167005899
			11'd1365: out = 32'b10000000000000000111110001101101; // input=-1.333984375, output=-0.972090844834
			11'd1366: out = 32'b10000000000000000111110010001011; // input=-1.337890625, output=-0.972999850858
			11'd1367: out = 32'b10000000000000000111110010101001; // input=-1.341796875, output=-0.973894010102
			11'd1368: out = 32'b10000000000000000111110011000101; // input=-1.345703125, output=-0.974773308922
			11'd1369: out = 32'b10000000000000000111110011100010; // input=-1.349609375, output=-0.9756377339
			11'd1370: out = 32'b10000000000000000111110011111110; // input=-1.353515625, output=-0.976487271847
			11'd1371: out = 32'b10000000000000000111110100011001; // input=-1.357421875, output=-0.977321909799
			11'd1372: out = 32'b10000000000000000111110100110100; // input=-1.361328125, output=-0.978141635021
			11'd1373: out = 32'b10000000000000000111110101001110; // input=-1.365234375, output=-0.978946435006
			11'd1374: out = 32'b10000000000000000111110101101000; // input=-1.369140625, output=-0.979736297472
			11'd1375: out = 32'b10000000000000000111110110000001; // input=-1.373046875, output=-0.980511210368
			11'd1376: out = 32'b10000000000000000111110110011010; // input=-1.376953125, output=-0.981271161869
			11'd1377: out = 32'b10000000000000000111110110110011; // input=-1.380859375, output=-0.98201614038
			11'd1378: out = 32'b10000000000000000111110111001011; // input=-1.384765625, output=-0.982746134532
			11'd1379: out = 32'b10000000000000000111110111100010; // input=-1.388671875, output=-0.983461133188
			11'd1380: out = 32'b10000000000000000111110111111001; // input=-1.392578125, output=-0.984161125436
			11'd1381: out = 32'b10000000000000000111111000001111; // input=-1.396484375, output=-0.984846100597
			11'd1382: out = 32'b10000000000000000111111000100101; // input=-1.400390625, output=-0.985516048218
			11'd1383: out = 32'b10000000000000000111111000111011; // input=-1.404296875, output=-0.986170958077
			11'd1384: out = 32'b10000000000000000111111001010000; // input=-1.408203125, output=-0.98681082018
			11'd1385: out = 32'b10000000000000000111111001100100; // input=-1.412109375, output=-0.987435624764
			11'd1386: out = 32'b10000000000000000111111001111000; // input=-1.416015625, output=-0.988045362295
			11'd1387: out = 32'b10000000000000000111111010001100; // input=-1.419921875, output=-0.98864002347
			11'd1388: out = 32'b10000000000000000111111010011111; // input=-1.423828125, output=-0.989219599214
			11'd1389: out = 32'b10000000000000000111111010110001; // input=-1.427734375, output=-0.989784080684
			11'd1390: out = 32'b10000000000000000111111011000011; // input=-1.431640625, output=-0.990333459267
			11'd1391: out = 32'b10000000000000000111111011010101; // input=-1.435546875, output=-0.99086772658
			11'd1392: out = 32'b10000000000000000111111011100110; // input=-1.439453125, output=-0.991386874471
			11'd1393: out = 32'b10000000000000000111111011110110; // input=-1.443359375, output=-0.991890895017
			11'd1394: out = 32'b10000000000000000111111100000110; // input=-1.447265625, output=-0.992379780529
			11'd1395: out = 32'b10000000000000000111111100010110; // input=-1.451171875, output=-0.992853523546
			11'd1396: out = 32'b10000000000000000111111100100101; // input=-1.455078125, output=-0.99331211684
			11'd1397: out = 32'b10000000000000000111111100110011; // input=-1.458984375, output=-0.993755553414
			11'd1398: out = 32'b10000000000000000111111101000001; // input=-1.462890625, output=-0.9941838265
			11'd1399: out = 32'b10000000000000000111111101001111; // input=-1.466796875, output=-0.994596929564
			11'd1400: out = 32'b10000000000000000111111101011100; // input=-1.470703125, output=-0.994994856303
			11'd1401: out = 32'b10000000000000000111111101101001; // input=-1.474609375, output=-0.995377600644
			11'd1402: out = 32'b10000000000000000111111101110101; // input=-1.478515625, output=-0.995745156748
			11'd1403: out = 32'b10000000000000000111111110000000; // input=-1.482421875, output=-0.996097519006
			11'd1404: out = 32'b10000000000000000111111110001011; // input=-1.486328125, output=-0.996434682041
			11'd1405: out = 32'b10000000000000000111111110010110; // input=-1.490234375, output=-0.996756640709
			11'd1406: out = 32'b10000000000000000111111110100000; // input=-1.494140625, output=-0.997063390097
			11'd1407: out = 32'b10000000000000000111111110101001; // input=-1.498046875, output=-0.997354925525
			11'd1408: out = 32'b10000000000000000111111110110010; // input=-1.501953125, output=-0.997631242543
			11'd1409: out = 32'b10000000000000000111111110111011; // input=-1.505859375, output=-0.997892336936
			11'd1410: out = 32'b10000000000000000111111111000011; // input=-1.509765625, output=-0.99813820472
			11'd1411: out = 32'b10000000000000000111111111001011; // input=-1.513671875, output=-0.998368842143
			11'd1412: out = 32'b10000000000000000111111111010010; // input=-1.517578125, output=-0.998584245685
			11'd1413: out = 32'b10000000000000000111111111011000; // input=-1.521484375, output=-0.998784412061
			11'd1414: out = 32'b10000000000000000111111111011110; // input=-1.525390625, output=-0.998969338215
			11'd1415: out = 32'b10000000000000000111111111100100; // input=-1.529296875, output=-0.999139021326
			11'd1416: out = 32'b10000000000000000111111111101001; // input=-1.533203125, output=-0.999293458805
			11'd1417: out = 32'b10000000000000000111111111101101; // input=-1.537109375, output=-0.999432648295
			11'd1418: out = 32'b10000000000000000111111111110001; // input=-1.541015625, output=-0.999556587673
			11'd1419: out = 32'b10000000000000000111111111110101; // input=-1.544921875, output=-0.999665275047
			11'd1420: out = 32'b10000000000000000111111111111000; // input=-1.548828125, output=-0.999758708759
			11'd1421: out = 32'b10000000000000000111111111111011; // input=-1.552734375, output=-0.999836887383
			11'd1422: out = 32'b10000000000000000111111111111101; // input=-1.556640625, output=-0.999899809726
			11'd1423: out = 32'b10000000000000000111111111111110; // input=-1.560546875, output=-0.999947474829
			11'd1424: out = 32'b10000000000000000111111111111111; // input=-1.564453125, output=-0.999979881963
			11'd1425: out = 32'b10000000000000000111111111111111; // input=-1.568359375, output=-0.999997030634
			11'd1426: out = 32'b10000000000000000111111111111111; // input=-1.572265625, output=-0.999998920582
			11'd1427: out = 32'b10000000000000000111111111111111; // input=-1.576171875, output=-0.999985551776
			11'd1428: out = 32'b10000000000000000111111111111111; // input=-1.580078125, output=-0.99995692442
			11'd1429: out = 32'b10000000000000000111111111111101; // input=-1.583984375, output=-0.999913038953
			11'd1430: out = 32'b10000000000000000111111111111011; // input=-1.587890625, output=-0.999853896042
			11'd1431: out = 32'b10000000000000000111111111111001; // input=-1.591796875, output=-0.999779496592
			11'd1432: out = 32'b10000000000000000111111111110110; // input=-1.595703125, output=-0.999689841736
			11'd1433: out = 32'b10000000000000000111111111110010; // input=-1.599609375, output=-0.999584932843
			11'd1434: out = 32'b10000000000000000111111111101110; // input=-1.603515625, output=-0.999464771514
			11'd1435: out = 32'b10000000000000000111111111101010; // input=-1.607421875, output=-0.999329359583
			11'd1436: out = 32'b10000000000000000111111111100101; // input=-1.611328125, output=-0.999178699114
			11'd1437: out = 32'b10000000000000000111111111100000; // input=-1.615234375, output=-0.999012792408
			11'd1438: out = 32'b10000000000000000111111111011010; // input=-1.619140625, output=-0.998831641997
			11'd1439: out = 32'b10000000000000000111111111010011; // input=-1.623046875, output=-0.998635250643
			11'd1440: out = 32'b10000000000000000111111111001100; // input=-1.626953125, output=-0.998423621343
			11'd1441: out = 32'b10000000000000000111111111000101; // input=-1.630859375, output=-0.998196757328
			11'd1442: out = 32'b10000000000000000111111110111101; // input=-1.634765625, output=-0.997954662059
			11'd1443: out = 32'b10000000000000000111111110110101; // input=-1.638671875, output=-0.997697339229
			11'd1444: out = 32'b10000000000000000111111110101100; // input=-1.642578125, output=-0.997424792765
			11'd1445: out = 32'b10000000000000000111111110100010; // input=-1.646484375, output=-0.997137026826
			11'd1446: out = 32'b10000000000000000111111110011000; // input=-1.650390625, output=-0.996834045803
			11'd1447: out = 32'b10000000000000000111111110001110; // input=-1.654296875, output=-0.996515854318
			11'd1448: out = 32'b10000000000000000111111110000011; // input=-1.658203125, output=-0.996182457228
			11'd1449: out = 32'b10000000000000000111111101110111; // input=-1.662109375, output=-0.995833859619
			11'd1450: out = 32'b10000000000000000111111101101100; // input=-1.666015625, output=-0.995470066811
			11'd1451: out = 32'b10000000000000000111111101011111; // input=-1.669921875, output=-0.995091084354
			11'd1452: out = 32'b10000000000000000111111101010010; // input=-1.673828125, output=-0.994696918032
			11'd1453: out = 32'b10000000000000000111111101000101; // input=-1.677734375, output=-0.994287573858
			11'd1454: out = 32'b10000000000000000111111100110111; // input=-1.681640625, output=-0.99386305808
			11'd1455: out = 32'b10000000000000000111111100101000; // input=-1.685546875, output=-0.993423377174
			11'd1456: out = 32'b10000000000000000111111100011010; // input=-1.689453125, output=-0.992968537849
			11'd1457: out = 32'b10000000000000000111111100001010; // input=-1.693359375, output=-0.992498547046
			11'd1458: out = 32'b10000000000000000111111011111010; // input=-1.697265625, output=-0.992013411937
			11'd1459: out = 32'b10000000000000000111111011101010; // input=-1.701171875, output=-0.991513139923
			11'd1460: out = 32'b10000000000000000111111011011001; // input=-1.705078125, output=-0.990997738639
			11'd1461: out = 32'b10000000000000000111111011001000; // input=-1.708984375, output=-0.990467215948
			11'd1462: out = 32'b10000000000000000111111010110110; // input=-1.712890625, output=-0.989921579947
			11'd1463: out = 32'b10000000000000000111111010100011; // input=-1.716796875, output=-0.98936083896
			11'd1464: out = 32'b10000000000000000111111010010001; // input=-1.720703125, output=-0.988785001544
			11'd1465: out = 32'b10000000000000000111111001111101; // input=-1.724609375, output=-0.988194076485
			11'd1466: out = 32'b10000000000000000111111001101001; // input=-1.728515625, output=-0.9875880728
			11'd1467: out = 32'b10000000000000000111111001010101; // input=-1.732421875, output=-0.986966999737
			11'd1468: out = 32'b10000000000000000111111001000000; // input=-1.736328125, output=-0.986330866772
			11'd1469: out = 32'b10000000000000000111111000101011; // input=-1.740234375, output=-0.98567968361
			11'd1470: out = 32'b10000000000000000111111000010101; // input=-1.744140625, output=-0.98501346019
			11'd1471: out = 32'b10000000000000000111110111111111; // input=-1.748046875, output=-0.984332206676
			11'd1472: out = 32'b10000000000000000111110111101000; // input=-1.751953125, output=-0.983635933464
			11'd1473: out = 32'b10000000000000000111110111010000; // input=-1.755859375, output=-0.982924651178
			11'd1474: out = 32'b10000000000000000111110110111001; // input=-1.759765625, output=-0.982198370671
			11'd1475: out = 32'b10000000000000000111110110100000; // input=-1.763671875, output=-0.981457103025
			11'd1476: out = 32'b10000000000000000111110110001000; // input=-1.767578125, output=-0.980700859551
			11'd1477: out = 32'b10000000000000000111110101101110; // input=-1.771484375, output=-0.979929651789
			11'd1478: out = 32'b10000000000000000111110101010101; // input=-1.775390625, output=-0.979143491506
			11'd1479: out = 32'b10000000000000000111110100111010; // input=-1.779296875, output=-0.978342390698
			11'd1480: out = 32'b10000000000000000111110100100000; // input=-1.783203125, output=-0.977526361588
			11'd1481: out = 32'b10000000000000000111110100000100; // input=-1.787109375, output=-0.976695416629
			11'd1482: out = 32'b10000000000000000111110011101001; // input=-1.791015625, output=-0.9758495685
			11'd1483: out = 32'b10000000000000000111110011001100; // input=-1.794921875, output=-0.974988830107
			11'd1484: out = 32'b10000000000000000111110010110000; // input=-1.798828125, output=-0.974113214584
			11'd1485: out = 32'b10000000000000000111110010010011; // input=-1.802734375, output=-0.973222735292
			11'd1486: out = 32'b10000000000000000111110001110101; // input=-1.806640625, output=-0.972317405818
			11'd1487: out = 32'b10000000000000000111110001010111; // input=-1.810546875, output=-0.971397239977
			11'd1488: out = 32'b10000000000000000111110000111000; // input=-1.814453125, output=-0.970462251809
			11'd1489: out = 32'b10000000000000000111110000011001; // input=-1.818359375, output=-0.969512455581
			11'd1490: out = 32'b10000000000000000111101111111001; // input=-1.822265625, output=-0.968547865786
			11'd1491: out = 32'b10000000000000000111101111011001; // input=-1.826171875, output=-0.967568497142
			11'd1492: out = 32'b10000000000000000111101110111001; // input=-1.830078125, output=-0.966574364594
			11'd1493: out = 32'b10000000000000000111101110011000; // input=-1.833984375, output=-0.96556548331
			11'd1494: out = 32'b10000000000000000111101101110110; // input=-1.837890625, output=-0.964541868684
			11'd1495: out = 32'b10000000000000000111101101010100; // input=-1.841796875, output=-0.963503536336
			11'd1496: out = 32'b10000000000000000111101100110010; // input=-1.845703125, output=-0.96245050211
			11'd1497: out = 32'b10000000000000000111101100001111; // input=-1.849609375, output=-0.961382782073
			11'd1498: out = 32'b10000000000000000111101011101011; // input=-1.853515625, output=-0.960300392518
			11'd1499: out = 32'b10000000000000000111101011000111; // input=-1.857421875, output=-0.95920334996
			11'd1500: out = 32'b10000000000000000111101010100011; // input=-1.861328125, output=-0.95809167114
			11'd1501: out = 32'b10000000000000000111101001111110; // input=-1.865234375, output=-0.956965373019
			11'd1502: out = 32'b10000000000000000111101001011000; // input=-1.869140625, output=-0.955824472784
			11'd1503: out = 32'b10000000000000000111101000110011; // input=-1.873046875, output=-0.954668987843
			11'd1504: out = 32'b10000000000000000111101000001100; // input=-1.876953125, output=-0.953498935829
			11'd1505: out = 32'b10000000000000000111100111100101; // input=-1.880859375, output=-0.952314334593
			11'd1506: out = 32'b10000000000000000111100110111110; // input=-1.884765625, output=-0.951115202213
			11'd1507: out = 32'b10000000000000000111100110010110; // input=-1.888671875, output=-0.949901556985
			11'd1508: out = 32'b10000000000000000111100101101110; // input=-1.892578125, output=-0.948673417428
			11'd1509: out = 32'b10000000000000000111100101000101; // input=-1.896484375, output=-0.947430802281
			11'd1510: out = 32'b10000000000000000111100100011100; // input=-1.900390625, output=-0.946173730507
			11'd1511: out = 32'b10000000000000000111100011110011; // input=-1.904296875, output=-0.944902221285
			11'd1512: out = 32'b10000000000000000111100011001000; // input=-1.908203125, output=-0.943616294018
			11'd1513: out = 32'b10000000000000000111100010011110; // input=-1.912109375, output=-0.942315968327
			11'd1514: out = 32'b10000000000000000111100001110011; // input=-1.916015625, output=-0.941001264054
			11'd1515: out = 32'b10000000000000000111100001000111; // input=-1.919921875, output=-0.939672201259
			11'd1516: out = 32'b10000000000000000111100000011011; // input=-1.923828125, output=-0.938328800223
			11'd1517: out = 32'b10000000000000000111011111101111; // input=-1.927734375, output=-0.936971081444
			11'd1518: out = 32'b10000000000000000111011111000010; // input=-1.931640625, output=-0.935599065638
			11'd1519: out = 32'b10000000000000000111011110010100; // input=-1.935546875, output=-0.934212773742
			11'd1520: out = 32'b10000000000000000111011101100110; // input=-1.939453125, output=-0.932812226909
			11'd1521: out = 32'b10000000000000000111011100111000; // input=-1.943359375, output=-0.931397446509
			11'd1522: out = 32'b10000000000000000111011100001001; // input=-1.947265625, output=-0.929968454129
			11'd1523: out = 32'b10000000000000000111011011011010; // input=-1.951171875, output=-0.928525271575
			11'd1524: out = 32'b10000000000000000111011010101010; // input=-1.955078125, output=-0.927067920868
			11'd1525: out = 32'b10000000000000000111011001111010; // input=-1.958984375, output=-0.925596424245
			11'd1526: out = 32'b10000000000000000111011001001001; // input=-1.962890625, output=-0.92411080416
			11'd1527: out = 32'b10000000000000000111011000011000; // input=-1.966796875, output=-0.92261108328
			11'd1528: out = 32'b10000000000000000111010111100111; // input=-1.970703125, output=-0.921097284491
			11'd1529: out = 32'b10000000000000000111010110110100; // input=-1.974609375, output=-0.91956943089
			11'd1530: out = 32'b10000000000000000111010110000010; // input=-1.978515625, output=-0.918027545791
			11'd1531: out = 32'b10000000000000000111010101001111; // input=-1.982421875, output=-0.916471652721
			11'd1532: out = 32'b10000000000000000111010100011100; // input=-1.986328125, output=-0.914901775422
			11'd1533: out = 32'b10000000000000000111010011101000; // input=-1.990234375, output=-0.913317937847
			11'd1534: out = 32'b10000000000000000111010010110011; // input=-1.994140625, output=-0.911720164164
			11'd1535: out = 32'b10000000000000000111010001111110; // input=-1.998046875, output=-0.910108478752
			11'd1536: out = 32'b10000000000000000111010001001001; // input=-2.001953125, output=-0.908482906206
			11'd1537: out = 32'b10000000000000000111010000010011; // input=-2.005859375, output=-0.906843471327
			11'd1538: out = 32'b10000000000000000111001111011101; // input=-2.009765625, output=-0.905190199134
			11'd1539: out = 32'b10000000000000000111001110100111; // input=-2.013671875, output=-0.903523114851
			11'd1540: out = 32'b10000000000000000111001101110000; // input=-2.017578125, output=-0.901842243918
			11'd1541: out = 32'b10000000000000000111001100111000; // input=-2.021484375, output=-0.900147611981
			11'd1542: out = 32'b10000000000000000111001100000000; // input=-2.025390625, output=-0.898439244899
			11'd1543: out = 32'b10000000000000000111001011001000; // input=-2.029296875, output=-0.89671716874
			11'd1544: out = 32'b10000000000000000111001010001111; // input=-2.033203125, output=-0.89498140978
			11'd1545: out = 32'b10000000000000000111001001010101; // input=-2.037109375, output=-0.893231994505
			11'd1546: out = 32'b10000000000000000111001000011100; // input=-2.041015625, output=-0.891468949608
			11'd1547: out = 32'b10000000000000000111000111100001; // input=-2.044921875, output=-0.889692301992
			11'd1548: out = 32'b10000000000000000111000110100111; // input=-2.048828125, output=-0.887902078767
			11'd1549: out = 32'b10000000000000000111000101101100; // input=-2.052734375, output=-0.886098307248
			11'd1550: out = 32'b10000000000000000111000100110000; // input=-2.056640625, output=-0.884281014959
			11'd1551: out = 32'b10000000000000000111000011110100; // input=-2.060546875, output=-0.882450229629
			11'd1552: out = 32'b10000000000000000111000010111000; // input=-2.064453125, output=-0.880605979195
			11'd1553: out = 32'b10000000000000000111000001111011; // input=-2.068359375, output=-0.878748291797
			11'd1554: out = 32'b10000000000000000111000000111110; // input=-2.072265625, output=-0.876877195782
			11'd1555: out = 32'b10000000000000000111000000000000; // input=-2.076171875, output=-0.874992719699
			11'd1556: out = 32'b10000000000000000110111111000010; // input=-2.080078125, output=-0.873094892304
			11'd1557: out = 32'b10000000000000000110111110000011; // input=-2.083984375, output=-0.871183742555
			11'd1558: out = 32'b10000000000000000110111101000100; // input=-2.087890625, output=-0.869259299614
			11'd1559: out = 32'b10000000000000000110111100000100; // input=-2.091796875, output=-0.867321592845
			11'd1560: out = 32'b10000000000000000110111011000100; // input=-2.095703125, output=-0.865370651816
			11'd1561: out = 32'b10000000000000000110111010000100; // input=-2.099609375, output=-0.863406506296
			11'd1562: out = 32'b10000000000000000110111001000011; // input=-2.103515625, output=-0.861429186254
			11'd1563: out = 32'b10000000000000000110111000000010; // input=-2.107421875, output=-0.859438721864
			11'd1564: out = 32'b10000000000000000110110111000000; // input=-2.111328125, output=-0.857435143495
			11'd1565: out = 32'b10000000000000000110110101111110; // input=-2.115234375, output=-0.855418481721
			11'd1566: out = 32'b10000000000000000110110100111100; // input=-2.119140625, output=-0.853388767314
			11'd1567: out = 32'b10000000000000000110110011111001; // input=-2.123046875, output=-0.851346031244
			11'd1568: out = 32'b10000000000000000110110010110110; // input=-2.126953125, output=-0.849290304681
			11'd1569: out = 32'b10000000000000000110110001110010; // input=-2.130859375, output=-0.847221618993
			11'd1570: out = 32'b10000000000000000110110000101110; // input=-2.134765625, output=-0.845140005746
			11'd1571: out = 32'b10000000000000000110101111101001; // input=-2.138671875, output=-0.843045496701
			11'd1572: out = 32'b10000000000000000110101110100100; // input=-2.142578125, output=-0.84093812382
			11'd1573: out = 32'b10000000000000000110101101011110; // input=-2.146484375, output=-0.838817919257
			11'd1574: out = 32'b10000000000000000110101100011000; // input=-2.150390625, output=-0.836684915366
			11'd1575: out = 32'b10000000000000000110101011010010; // input=-2.154296875, output=-0.834539144691
			11'd1576: out = 32'b10000000000000000110101010001011; // input=-2.158203125, output=-0.832380639976
			11'd1577: out = 32'b10000000000000000110101001000100; // input=-2.162109375, output=-0.830209434157
			11'd1578: out = 32'b10000000000000000110100111111101; // input=-2.166015625, output=-0.828025560363
			11'd1579: out = 32'b10000000000000000110100110110101; // input=-2.169921875, output=-0.825829051918
			11'd1580: out = 32'b10000000000000000110100101101100; // input=-2.173828125, output=-0.823619942338
			11'd1581: out = 32'b10000000000000000110100100100100; // input=-2.177734375, output=-0.82139826533
			11'd1582: out = 32'b10000000000000000110100011011010; // input=-2.181640625, output=-0.819164054796
			11'd1583: out = 32'b10000000000000000110100010010001; // input=-2.185546875, output=-0.816917344826
			11'd1584: out = 32'b10000000000000000110100001000111; // input=-2.189453125, output=-0.814658169702
			11'd1585: out = 32'b10000000000000000110011111111100; // input=-2.193359375, output=-0.812386563897
			11'd1586: out = 32'b10000000000000000110011110110001; // input=-2.197265625, output=-0.810102562073
			11'd1587: out = 32'b10000000000000000110011101100110; // input=-2.201171875, output=-0.80780619908
			11'd1588: out = 32'b10000000000000000110011100011011; // input=-2.205078125, output=-0.805497509959
			11'd1589: out = 32'b10000000000000000110011011001110; // input=-2.208984375, output=-0.803176529936
			11'd1590: out = 32'b10000000000000000110011010000010; // input=-2.212890625, output=-0.800843294428
			11'd1591: out = 32'b10000000000000000110011000110101; // input=-2.216796875, output=-0.798497839037
			11'd1592: out = 32'b10000000000000000110010111101000; // input=-2.220703125, output=-0.796140199551
			11'd1593: out = 32'b10000000000000000110010110011010; // input=-2.224609375, output=-0.793770411945
			11'd1594: out = 32'b10000000000000000110010101001100; // input=-2.228515625, output=-0.791388512379
			11'd1595: out = 32'b10000000000000000110010011111110; // input=-2.232421875, output=-0.788994537198
			11'd1596: out = 32'b10000000000000000110010010101111; // input=-2.236328125, output=-0.786588522931
			11'd1597: out = 32'b10000000000000000110010001100000; // input=-2.240234375, output=-0.784170506291
			11'd1598: out = 32'b10000000000000000110010000010000; // input=-2.244140625, output=-0.781740524174
			11'd1599: out = 32'b10000000000000000110001111000000; // input=-2.248046875, output=-0.779298613658
			11'd1600: out = 32'b10000000000000000110001101110000; // input=-2.251953125, output=-0.776844812005
			11'd1601: out = 32'b10000000000000000110001100011111; // input=-2.255859375, output=-0.774379156655
			11'd1602: out = 32'b10000000000000000110001011001110; // input=-2.259765625, output=-0.771901685232
			11'd1603: out = 32'b10000000000000000110001001111100; // input=-2.263671875, output=-0.769412435539
			11'd1604: out = 32'b10000000000000000110001000101010; // input=-2.267578125, output=-0.766911445559
			11'd1605: out = 32'b10000000000000000110000111011000; // input=-2.271484375, output=-0.764398753454
			11'd1606: out = 32'b10000000000000000110000110000101; // input=-2.275390625, output=-0.761874397564
			11'd1607: out = 32'b10000000000000000110000100110010; // input=-2.279296875, output=-0.759338416409
			11'd1608: out = 32'b10000000000000000110000011011111; // input=-2.283203125, output=-0.756790848683
			11'd1609: out = 32'b10000000000000000110000010001011; // input=-2.287109375, output=-0.75423173326
			11'd1610: out = 32'b10000000000000000110000000110110; // input=-2.291015625, output=-0.751661109189
			11'd1611: out = 32'b10000000000000000101111111100010; // input=-2.294921875, output=-0.749079015694
			11'd1612: out = 32'b10000000000000000101111110001101; // input=-2.298828125, output=-0.746485492175
			11'd1613: out = 32'b10000000000000000101111100110111; // input=-2.302734375, output=-0.743880578206
			11'd1614: out = 32'b10000000000000000101111011100010; // input=-2.306640625, output=-0.741264313535
			11'd1615: out = 32'b10000000000000000101111010001100; // input=-2.310546875, output=-0.738636738082
			11'd1616: out = 32'b10000000000000000101111000110101; // input=-2.314453125, output=-0.735997891941
			11'd1617: out = 32'b10000000000000000101110111011110; // input=-2.318359375, output=-0.733347815378
			11'd1618: out = 32'b10000000000000000101110110000111; // input=-2.322265625, output=-0.730686548829
			11'd1619: out = 32'b10000000000000000101110100110000; // input=-2.326171875, output=-0.728014132903
			11'd1620: out = 32'b10000000000000000101110011011000; // input=-2.330078125, output=-0.725330608377
			11'd1621: out = 32'b10000000000000000101110001111111; // input=-2.333984375, output=-0.722636016198
			11'd1622: out = 32'b10000000000000000101110000100111; // input=-2.337890625, output=-0.719930397482
			11'd1623: out = 32'b10000000000000000101101111001110; // input=-2.341796875, output=-0.717213793515
			11'd1624: out = 32'b10000000000000000101101101110100; // input=-2.345703125, output=-0.714486245747
			11'd1625: out = 32'b10000000000000000101101100011011; // input=-2.349609375, output=-0.711747795798
			11'd1626: out = 32'b10000000000000000101101011000000; // input=-2.353515625, output=-0.708998485454
			11'd1627: out = 32'b10000000000000000101101001100110; // input=-2.357421875, output=-0.706238356665
			11'd1628: out = 32'b10000000000000000101101000001011; // input=-2.361328125, output=-0.703467451548
			11'd1629: out = 32'b10000000000000000101100110110000; // input=-2.365234375, output=-0.700685812383
			11'd1630: out = 32'b10000000000000000101100101010101; // input=-2.369140625, output=-0.697893481614
			11'd1631: out = 32'b10000000000000000101100011111001; // input=-2.373046875, output=-0.69509050185
			11'd1632: out = 32'b10000000000000000101100010011101; // input=-2.376953125, output=-0.692276915859
			11'd1633: out = 32'b10000000000000000101100001000000; // input=-2.380859375, output=-0.689452766575
			11'd1634: out = 32'b10000000000000000101011111100011; // input=-2.384765625, output=-0.68661809709
			11'd1635: out = 32'b10000000000000000101011110000110; // input=-2.388671875, output=-0.683772950657
			11'd1636: out = 32'b10000000000000000101011100101000; // input=-2.392578125, output=-0.680917370691
			11'd1637: out = 32'b10000000000000000101011011001010; // input=-2.396484375, output=-0.678051400763
			11'd1638: out = 32'b10000000000000000101011001101100; // input=-2.400390625, output=-0.675175084605
			11'd1639: out = 32'b10000000000000000101011000001110; // input=-2.404296875, output=-0.672288466105
			11'd1640: out = 32'b10000000000000000101010110101111; // input=-2.408203125, output=-0.669391589311
			11'd1641: out = 32'b10000000000000000101010101001111; // input=-2.412109375, output=-0.666484498425
			11'd1642: out = 32'b10000000000000000101010011110000; // input=-2.416015625, output=-0.663567237806
			11'd1643: out = 32'b10000000000000000101010010010000; // input=-2.419921875, output=-0.660639851967
			11'd1644: out = 32'b10000000000000000101010000110000; // input=-2.423828125, output=-0.657702385576
			11'd1645: out = 32'b10000000000000000101001111001111; // input=-2.427734375, output=-0.654754883457
			11'd1646: out = 32'b10000000000000000101001101101110; // input=-2.431640625, output=-0.651797390583
			11'd1647: out = 32'b10000000000000000101001100001101; // input=-2.435546875, output=-0.648829952083
			11'd1648: out = 32'b10000000000000000101001010101011; // input=-2.439453125, output=-0.645852613236
			11'd1649: out = 32'b10000000000000000101001001001001; // input=-2.443359375, output=-0.642865419473
			11'd1650: out = 32'b10000000000000000101000111100111; // input=-2.447265625, output=-0.639868416375
			11'd1651: out = 32'b10000000000000000101000110000101; // input=-2.451171875, output=-0.636861649672
			11'd1652: out = 32'b10000000000000000101000100100010; // input=-2.455078125, output=-0.633845165244
			11'd1653: out = 32'b10000000000000000101000010111111; // input=-2.458984375, output=-0.630819009118
			11'd1654: out = 32'b10000000000000000101000001011011; // input=-2.462890625, output=-0.62778322747
			11'd1655: out = 32'b10000000000000000100111111110111; // input=-2.466796875, output=-0.624737866623
			11'd1656: out = 32'b10000000000000000100111110010011; // input=-2.470703125, output=-0.621682973045
			11'd1657: out = 32'b10000000000000000100111100101111; // input=-2.474609375, output=-0.618618593349
			11'd1658: out = 32'b10000000000000000100111011001010; // input=-2.478515625, output=-0.615544774295
			11'd1659: out = 32'b10000000000000000100111001100101; // input=-2.482421875, output=-0.612461562784
			11'd1660: out = 32'b10000000000000000100111000000000; // input=-2.486328125, output=-0.609369005864
			11'd1661: out = 32'b10000000000000000100110110011010; // input=-2.490234375, output=-0.606267150722
			11'd1662: out = 32'b10000000000000000100110100110100; // input=-2.494140625, output=-0.60315604469
			11'd1663: out = 32'b10000000000000000100110011001110; // input=-2.498046875, output=-0.600035735239
			11'd1664: out = 32'b10000000000000000100110001100111; // input=-2.501953125, output=-0.59690626998
			11'd1665: out = 32'b10000000000000000100110000000001; // input=-2.505859375, output=-0.593767696666
			11'd1666: out = 32'b10000000000000000100101110011001; // input=-2.509765625, output=-0.590620063188
			11'd1667: out = 32'b10000000000000000100101100110010; // input=-2.513671875, output=-0.587463417574
			11'd1668: out = 32'b10000000000000000100101011001010; // input=-2.517578125, output=-0.584297807991
			11'd1669: out = 32'b10000000000000000100101001100010; // input=-2.521484375, output=-0.581123282743
			11'd1670: out = 32'b10000000000000000100100111111010; // input=-2.525390625, output=-0.577939890268
			11'd1671: out = 32'b10000000000000000100100110010001; // input=-2.529296875, output=-0.574747679141
			11'd1672: out = 32'b10000000000000000100100100101000; // input=-2.533203125, output=-0.571546698072
			11'd1673: out = 32'b10000000000000000100100010111111; // input=-2.537109375, output=-0.568336995904
			11'd1674: out = 32'b10000000000000000100100001010110; // input=-2.541015625, output=-0.565118621612
			11'd1675: out = 32'b10000000000000000100011111101100; // input=-2.544921875, output=-0.561891624306
			11'd1676: out = 32'b10000000000000000100011110000010; // input=-2.548828125, output=-0.558656053224
			11'd1677: out = 32'b10000000000000000100011100011000; // input=-2.552734375, output=-0.555411957739
			11'd1678: out = 32'b10000000000000000100011010101101; // input=-2.556640625, output=-0.55215938735
			11'd1679: out = 32'b10000000000000000100011001000010; // input=-2.560546875, output=-0.548898391689
			11'd1680: out = 32'b10000000000000000100010111010111; // input=-2.564453125, output=-0.545629020513
			11'd1681: out = 32'b10000000000000000100010101101100; // input=-2.568359375, output=-0.54235132371
			11'd1682: out = 32'b10000000000000000100010100000000; // input=-2.572265625, output=-0.539065351293
			11'd1683: out = 32'b10000000000000000100010010010100; // input=-2.576171875, output=-0.535771153402
			11'd1684: out = 32'b10000000000000000100010000101000; // input=-2.580078125, output=-0.532468780302
			11'd1685: out = 32'b10000000000000000100001110111011; // input=-2.583984375, output=-0.529158282384
			11'd1686: out = 32'b10000000000000000100001101001111; // input=-2.587890625, output=-0.525839710162
			11'd1687: out = 32'b10000000000000000100001011100010; // input=-2.591796875, output=-0.522513114272
			11'd1688: out = 32'b10000000000000000100001001110100; // input=-2.595703125, output=-0.519178545475
			11'd1689: out = 32'b10000000000000000100001000000111; // input=-2.599609375, output=-0.515836054653
			11'd1690: out = 32'b10000000000000000100000110011001; // input=-2.603515625, output=-0.512485692806
			11'd1691: out = 32'b10000000000000000100000100101011; // input=-2.607421875, output=-0.509127511059
			11'd1692: out = 32'b10000000000000000100000010111101; // input=-2.611328125, output=-0.505761560652
			11'd1693: out = 32'b10000000000000000100000001001110; // input=-2.615234375, output=-0.502387892946
			11'd1694: out = 32'b10000000000000000011111111011111; // input=-2.619140625, output=-0.499006559419
			11'd1695: out = 32'b10000000000000000011111101110000; // input=-2.623046875, output=-0.495617611666
			11'd1696: out = 32'b10000000000000000011111100000001; // input=-2.626953125, output=-0.492221101398
			11'd1697: out = 32'b10000000000000000011111010010010; // input=-2.630859375, output=-0.488817080442
			11'd1698: out = 32'b10000000000000000011111000100010; // input=-2.634765625, output=-0.485405600738
			11'd1699: out = 32'b10000000000000000011110110110010; // input=-2.638671875, output=-0.481986714342
			11'd1700: out = 32'b10000000000000000011110101000001; // input=-2.642578125, output=-0.478560473421
			11'd1701: out = 32'b10000000000000000011110011010001; // input=-2.646484375, output=-0.475126930257
			11'd1702: out = 32'b10000000000000000011110001100000; // input=-2.650390625, output=-0.47168613724
			11'd1703: out = 32'b10000000000000000011101111101111; // input=-2.654296875, output=-0.468238146873
			11'd1704: out = 32'b10000000000000000011101101111110; // input=-2.658203125, output=-0.464783011769
			11'd1705: out = 32'b10000000000000000011101100001101; // input=-2.662109375, output=-0.461320784647
			11'd1706: out = 32'b10000000000000000011101010011011; // input=-2.666015625, output=-0.457851518337
			11'd1707: out = 32'b10000000000000000011101000101001; // input=-2.669921875, output=-0.454375265777
			11'd1708: out = 32'b10000000000000000011100110110111; // input=-2.673828125, output=-0.450892080009
			11'd1709: out = 32'b10000000000000000011100101000100; // input=-2.677734375, output=-0.447402014183
			11'd1710: out = 32'b10000000000000000011100011010010; // input=-2.681640625, output=-0.443905121553
			11'd1711: out = 32'b10000000000000000011100001011111; // input=-2.685546875, output=-0.440401455476
			11'd1712: out = 32'b10000000000000000011011111101100; // input=-2.689453125, output=-0.436891069416
			11'd1713: out = 32'b10000000000000000011011101111001; // input=-2.693359375, output=-0.433374016935
			11'd1714: out = 32'b10000000000000000011011100000101; // input=-2.697265625, output=-0.429850351699
			11'd1715: out = 32'b10000000000000000011011010010010; // input=-2.701171875, output=-0.426320127476
			11'd1716: out = 32'b10000000000000000011011000011110; // input=-2.705078125, output=-0.422783398133
			11'd1717: out = 32'b10000000000000000011010110101010; // input=-2.708984375, output=-0.419240217635
			11'd1718: out = 32'b10000000000000000011010100110101; // input=-2.712890625, output=-0.415690640047
			11'd1719: out = 32'b10000000000000000011010011000001; // input=-2.716796875, output=-0.412134719532
			11'd1720: out = 32'b10000000000000000011010001001100; // input=-2.720703125, output=-0.408572510347
			11'd1721: out = 32'b10000000000000000011001111010111; // input=-2.724609375, output=-0.405004066849
			11'd1722: out = 32'b10000000000000000011001101100010; // input=-2.728515625, output=-0.401429443487
			11'd1723: out = 32'b10000000000000000011001011101101; // input=-2.732421875, output=-0.397848694806
			11'd1724: out = 32'b10000000000000000011001001110111; // input=-2.736328125, output=-0.394261875443
			11'd1725: out = 32'b10000000000000000011001000000001; // input=-2.740234375, output=-0.390669040129
			11'd1726: out = 32'b10000000000000000011000110001100; // input=-2.744140625, output=-0.387070243686
			11'd1727: out = 32'b10000000000000000011000100010101; // input=-2.748046875, output=-0.383465541027
			11'd1728: out = 32'b10000000000000000011000010011111; // input=-2.751953125, output=-0.379854987156
			11'd1729: out = 32'b10000000000000000011000000101001; // input=-2.755859375, output=-0.376238637166
			11'd1730: out = 32'b10000000000000000010111110110010; // input=-2.759765625, output=-0.372616546236
			11'd1731: out = 32'b10000000000000000010111100111011; // input=-2.763671875, output=-0.368988769637
			11'd1732: out = 32'b10000000000000000010111011000100; // input=-2.767578125, output=-0.365355362723
			11'd1733: out = 32'b10000000000000000010111001001101; // input=-2.771484375, output=-0.361716380935
			11'd1734: out = 32'b10000000000000000010110111010101; // input=-2.775390625, output=-0.358071879801
			11'd1735: out = 32'b10000000000000000010110101011110; // input=-2.779296875, output=-0.35442191493
			11'd1736: out = 32'b10000000000000000010110011100110; // input=-2.783203125, output=-0.350766542017
			11'd1737: out = 32'b10000000000000000010110001101110; // input=-2.787109375, output=-0.347105816838
			11'd1738: out = 32'b10000000000000000010101111110110; // input=-2.791015625, output=-0.343439795251
			11'd1739: out = 32'b10000000000000000010101101111110; // input=-2.794921875, output=-0.339768533196
			11'd1740: out = 32'b10000000000000000010101100000101; // input=-2.798828125, output=-0.336092086691
			11'd1741: out = 32'b10000000000000000010101010001100; // input=-2.802734375, output=-0.332410511834
			11'd1742: out = 32'b10000000000000000010101000010100; // input=-2.806640625, output=-0.328723864801
			11'd1743: out = 32'b10000000000000000010100110011011; // input=-2.810546875, output=-0.325032201847
			11'd1744: out = 32'b10000000000000000010100100100010; // input=-2.814453125, output=-0.321335579302
			11'd1745: out = 32'b10000000000000000010100010101000; // input=-2.818359375, output=-0.31763405357
			11'd1746: out = 32'b10000000000000000010100000101111; // input=-2.822265625, output=-0.313927681134
			11'd1747: out = 32'b10000000000000000010011110110101; // input=-2.826171875, output=-0.310216518548
			11'd1748: out = 32'b10000000000000000010011100111011; // input=-2.830078125, output=-0.306500622439
			11'd1749: out = 32'b10000000000000000010011011000001; // input=-2.833984375, output=-0.302780049508
			11'd1750: out = 32'b10000000000000000010011001000111; // input=-2.837890625, output=-0.299054856526
			11'd1751: out = 32'b10000000000000000010010111001101; // input=-2.841796875, output=-0.295325100335
			11'd1752: out = 32'b10000000000000000010010101010011; // input=-2.845703125, output=-0.291590837846
			11'd1753: out = 32'b10000000000000000010010011011000; // input=-2.849609375, output=-0.28785212604
			11'd1754: out = 32'b10000000000000000010010001011110; // input=-2.853515625, output=-0.284109021964
			11'd1755: out = 32'b10000000000000000010001111100011; // input=-2.857421875, output=-0.280361582734
			11'd1756: out = 32'b10000000000000000010001101101000; // input=-2.861328125, output=-0.276609865532
			11'd1757: out = 32'b10000000000000000010001011101101; // input=-2.865234375, output=-0.272853927603
			11'd1758: out = 32'b10000000000000000010001001110010; // input=-2.869140625, output=-0.269093826259
			11'd1759: out = 32'b10000000000000000010000111110110; // input=-2.873046875, output=-0.265329618874
			11'd1760: out = 32'b10000000000000000010000101111011; // input=-2.876953125, output=-0.261561362886
			11'd1761: out = 32'b10000000000000000010000011111111; // input=-2.880859375, output=-0.257789115793
			11'd1762: out = 32'b10000000000000000010000010000011; // input=-2.884765625, output=-0.254012935156
			11'd1763: out = 32'b10000000000000000010000000001000; // input=-2.888671875, output=-0.250232878593
			11'd1764: out = 32'b10000000000000000001111110001100; // input=-2.892578125, output=-0.246449003785
			11'd1765: out = 32'b10000000000000000001111100010000; // input=-2.896484375, output=-0.242661368468
			11'd1766: out = 32'b10000000000000000001111010010011; // input=-2.900390625, output=-0.238870030437
			11'd1767: out = 32'b10000000000000000001111000010111; // input=-2.904296875, output=-0.235075047543
			11'd1768: out = 32'b10000000000000000001110110011010; // input=-2.908203125, output=-0.231276477694
			11'd1769: out = 32'b10000000000000000001110100011110; // input=-2.912109375, output=-0.22747437885
			11'd1770: out = 32'b10000000000000000001110010100001; // input=-2.916015625, output=-0.223668809027
			11'd1771: out = 32'b10000000000000000001110000100100; // input=-2.919921875, output=-0.219859826292
			11'd1772: out = 32'b10000000000000000001101110100111; // input=-2.923828125, output=-0.216047488768
			11'd1773: out = 32'b10000000000000000001101100101010; // input=-2.927734375, output=-0.212231854624
			11'd1774: out = 32'b10000000000000000001101010101101; // input=-2.931640625, output=-0.208412982084
			11'd1775: out = 32'b10000000000000000001101000110000; // input=-2.935546875, output=-0.204590929418
			11'd1776: out = 32'b10000000000000000001100110110011; // input=-2.939453125, output=-0.200765754946
			11'd1777: out = 32'b10000000000000000001100100110101; // input=-2.943359375, output=-0.196937517036
			11'd1778: out = 32'b10000000000000000001100010111000; // input=-2.947265625, output=-0.193106274101
			11'd1779: out = 32'b10000000000000000001100000111010; // input=-2.951171875, output=-0.189272084602
			11'd1780: out = 32'b10000000000000000001011110111100; // input=-2.955078125, output=-0.185435007044
			11'd1781: out = 32'b10000000000000000001011100111111; // input=-2.958984375, output=-0.181595099977
			11'd1782: out = 32'b10000000000000000001011011000001; // input=-2.962890625, output=-0.177752421991
			11'd1783: out = 32'b10000000000000000001011001000011; // input=-2.966796875, output=-0.173907031722
			11'd1784: out = 32'b10000000000000000001010111000100; // input=-2.970703125, output=-0.170058987846
			11'd1785: out = 32'b10000000000000000001010101000110; // input=-2.974609375, output=-0.166208349078
			11'd1786: out = 32'b10000000000000000001010011001000; // input=-2.978515625, output=-0.162355174176
			11'd1787: out = 32'b10000000000000000001010001001010; // input=-2.982421875, output=-0.158499521934
			11'd1788: out = 32'b10000000000000000001001111001011; // input=-2.986328125, output=-0.154641451184
			11'd1789: out = 32'b10000000000000000001001101001101; // input=-2.990234375, output=-0.150781020795
			11'd1790: out = 32'b10000000000000000001001011001110; // input=-2.994140625, output=-0.146918289674
			11'd1791: out = 32'b10000000000000000001001001010000; // input=-2.998046875, output=-0.14305331676
			11'd1792: out = 32'b10000000000000000001000111010001; // input=-3.001953125, output=-0.139186161029
			11'd1793: out = 32'b10000000000000000001000101010010; // input=-3.005859375, output=-0.135316881489
			11'd1794: out = 32'b10000000000000000001000011010011; // input=-3.009765625, output=-0.131445537179
			11'd1795: out = 32'b10000000000000000001000001010100; // input=-3.013671875, output=-0.127572187172
			11'd1796: out = 32'b10000000000000000000111111010101; // input=-3.017578125, output=-0.12369689057
			11'd1797: out = 32'b10000000000000000000111101010110; // input=-3.021484375, output=-0.119819706506
			11'd1798: out = 32'b10000000000000000000111011010111; // input=-3.025390625, output=-0.115940694141
			11'd1799: out = 32'b10000000000000000000111001011000; // input=-3.029296875, output=-0.112059912663
			11'd1800: out = 32'b10000000000000000000110111011001; // input=-3.033203125, output=-0.108177421289
			11'd1801: out = 32'b10000000000000000000110101011001; // input=-3.037109375, output=-0.10429327926
			11'd1802: out = 32'b10000000000000000000110011011010; // input=-3.041015625, output=-0.100407545845
			11'd1803: out = 32'b10000000000000000000110001011011; // input=-3.044921875, output=-0.0965202803338
			11'd1804: out = 32'b10000000000000000000101111011011; // input=-3.048828125, output=-0.0926315420419
			11'd1805: out = 32'b10000000000000000000101101011100; // input=-3.052734375, output=-0.0887413903066
			11'd1806: out = 32'b10000000000000000000101011011100; // input=-3.056640625, output=-0.0848498844869
			11'd1807: out = 32'b10000000000000000000101001011101; // input=-3.060546875, output=-0.0809570839624
			11'd1808: out = 32'b10000000000000000000100111011101; // input=-3.064453125, output=-0.0770630481324
			11'd1809: out = 32'b10000000000000000000100101011110; // input=-3.068359375, output=-0.0731678364151
			11'd1810: out = 32'b10000000000000000000100011011110; // input=-3.072265625, output=-0.0692715082466
			11'd1811: out = 32'b10000000000000000000100001011110; // input=-3.076171875, output=-0.0653741230801
			11'd1812: out = 32'b10000000000000000000011111011110; // input=-3.080078125, output=-0.061475740385
			11'd1813: out = 32'b10000000000000000000011101011111; // input=-3.083984375, output=-0.0575764196456
			11'd1814: out = 32'b10000000000000000000011011011111; // input=-3.087890625, output=-0.053676220361
			11'd1815: out = 32'b10000000000000000000011001011111; // input=-3.091796875, output=-0.0497752020432
			11'd1816: out = 32'b10000000000000000000010111011111; // input=-3.095703125, output=-0.0458734242172
			11'd1817: out = 32'b10000000000000000000010101011111; // input=-3.099609375, output=-0.0419709464191
			11'd1818: out = 32'b10000000000000000000010011011111; // input=-3.103515625, output=-0.038067828196
			11'd1819: out = 32'b10000000000000000000010001011111; // input=-3.107421875, output=-0.0341641291047
			11'd1820: out = 32'b10000000000000000000001111100000; // input=-3.111328125, output=-0.0302599087108
			11'd1821: out = 32'b10000000000000000000001101100000; // input=-3.115234375, output=-0.0263552265879
			11'd1822: out = 32'b10000000000000000000001011100000; // input=-3.119140625, output=-0.0224501423167
			11'd1823: out = 32'b10000000000000000000001001100000; // input=-3.123046875, output=-0.018544715484
			11'd1824: out = 32'b10000000000000000000000111100000; // input=-3.126953125, output=-0.0146390056817
			11'd1825: out = 32'b10000000000000000000000101100000; // input=-3.130859375, output=-0.0107330725062
			11'd1826: out = 32'b10000000000000000000000011100000; // input=-3.134765625, output=-0.0068269755572
			11'd1827: out = 32'b10000000000000000000000001100000; // input=-3.138671875, output=-0.00292077443696
			11'd1828: out = 32'b00000000000000000000000000100000; // input=-3.142578125, output=0.000985471250699
			11'd1829: out = 32'b00000000000000000000000010100000; // input=-3.146484375, output=0.00489170190128
			11'd1830: out = 32'b00000000000000000000000100100000; // input=-3.150390625, output=0.00879785791051
			11'd1831: out = 32'b00000000000000000000000110100000; // input=-3.154296875, output=0.0127038796752
			11'd1832: out = 32'b00000000000000000000001000100000; // input=-3.158203125, output=0.0166097075944
			11'd1833: out = 32'b00000000000000000000001010100000; // input=-3.162109375, output=0.0205152820699
			11'd1834: out = 32'b00000000000000000000001100100000; // input=-3.166015625, output=0.0244205435074
			11'd1835: out = 32'b00000000000000000000001110100000; // input=-3.169921875, output=0.0283254323174
			11'd1836: out = 32'b00000000000000000000010000100000; // input=-3.173828125, output=0.0322298889162
			11'd1837: out = 32'b00000000000000000000010010100000; // input=-3.177734375, output=0.0361338537266
			11'd1838: out = 32'b00000000000000000000010100100000; // input=-3.181640625, output=0.0400372671788
			11'd1839: out = 32'b00000000000000000000010110100000; // input=-3.185546875, output=0.0439400697116
			11'd1840: out = 32'b00000000000000000000011000100000; // input=-3.189453125, output=0.0478422017729
			11'd1841: out = 32'b00000000000000000000011010100000; // input=-3.193359375, output=0.0517436038212
			11'd1842: out = 32'b00000000000000000000011100011111; // input=-3.197265625, output=0.0556442163256
			11'd1843: out = 32'b00000000000000000000011110011111; // input=-3.201171875, output=0.0595439797679
			11'd1844: out = 32'b00000000000000000000100000011111; // input=-3.205078125, output=0.0634428346422
			11'd1845: out = 32'b00000000000000000000100010011111; // input=-3.208984375, output=0.0673407214569
			11'd1846: out = 32'b00000000000000000000100100011110; // input=-3.212890625, output=0.0712375807351
			11'd1847: out = 32'b00000000000000000000100110011110; // input=-3.216796875, output=0.0751333530155
			11'd1848: out = 32'b00000000000000000000101000011110; // input=-3.220703125, output=0.0790279788533
			11'd1849: out = 32'b00000000000000000000101010011101; // input=-3.224609375, output=0.0829213988214
			11'd1850: out = 32'b00000000000000000000101100011101; // input=-3.228515625, output=0.086813553511
			11'd1851: out = 32'b00000000000000000000101110011100; // input=-3.232421875, output=0.0907043835325
			11'd1852: out = 32'b00000000000000000000110000011100; // input=-3.236328125, output=0.0945938295168
			11'd1853: out = 32'b00000000000000000000110010011011; // input=-3.240234375, output=0.0984818321156
			11'd1854: out = 32'b00000000000000000000110100011010; // input=-3.244140625, output=0.102368332003
			11'd1855: out = 32'b00000000000000000000110110011010; // input=-3.248046875, output=0.106253269875
			11'd1856: out = 32'b00000000000000000000111000011001; // input=-3.251953125, output=0.110136586453
			11'd1857: out = 32'b00000000000000000000111010011000; // input=-3.255859375, output=0.114018222483
			11'd1858: out = 32'b00000000000000000000111100010111; // input=-3.259765625, output=0.117898118735
			11'd1859: out = 32'b00000000000000000000111110010110; // input=-3.263671875, output=0.121776216006
			11'd1860: out = 32'b00000000000000000001000000010101; // input=-3.267578125, output=0.125652455122
			11'd1861: out = 32'b00000000000000000001000010010100; // input=-3.271484375, output=0.129526776936
			11'd1862: out = 32'b00000000000000000001000100010011; // input=-3.275390625, output=0.133399122331
			11'd1863: out = 32'b00000000000000000001000110010010; // input=-3.279296875, output=0.13726943222
			11'd1864: out = 32'b00000000000000000001001000010001; // input=-3.283203125, output=0.141137647546
			11'd1865: out = 32'b00000000000000000001001010001111; // input=-3.287109375, output=0.145003709285
			11'd1866: out = 32'b00000000000000000001001100001110; // input=-3.291015625, output=0.148867558446
			11'd1867: out = 32'b00000000000000000001001110001101; // input=-3.294921875, output=0.152729136071
			11'd1868: out = 32'b00000000000000000001010000001011; // input=-3.298828125, output=0.156588383237
			11'd1869: out = 32'b00000000000000000001010010001001; // input=-3.302734375, output=0.160445241058
			11'd1870: out = 32'b00000000000000000001010100001000; // input=-3.306640625, output=0.164299650681
			11'd1871: out = 32'b00000000000000000001010110000110; // input=-3.310546875, output=0.168151553294
			11'd1872: out = 32'b00000000000000000001011000000100; // input=-3.314453125, output=0.172000890121
			11'd1873: out = 32'b00000000000000000001011010000010; // input=-3.318359375, output=0.175847602426
			11'd1874: out = 32'b00000000000000000001011100000000; // input=-3.322265625, output=0.179691631513
			11'd1875: out = 32'b00000000000000000001011101111110; // input=-3.326171875, output=0.183532918727
			11'd1876: out = 32'b00000000000000000001011111111100; // input=-3.330078125, output=0.187371405454
			11'd1877: out = 32'b00000000000000000001100001111001; // input=-3.333984375, output=0.191207033124
			11'd1878: out = 32'b00000000000000000001100011110111; // input=-3.337890625, output=0.19503974321
			11'd1879: out = 32'b00000000000000000001100101110101; // input=-3.341796875, output=0.198869477229
			11'd1880: out = 32'b00000000000000000001100111110010; // input=-3.345703125, output=0.202696176745
			11'd1881: out = 32'b00000000000000000001101001101111; // input=-3.349609375, output=0.206519783367
			11'd1882: out = 32'b00000000000000000001101011101100; // input=-3.353515625, output=0.210340238751
			11'd1883: out = 32'b00000000000000000001101101101010; // input=-3.357421875, output=0.214157484602
			11'd1884: out = 32'b00000000000000000001101111100110; // input=-3.361328125, output=0.217971462672
			11'd1885: out = 32'b00000000000000000001110001100011; // input=-3.365234375, output=0.221782114767
			11'd1886: out = 32'b00000000000000000001110011100000; // input=-3.369140625, output=0.225589382739
			11'd1887: out = 32'b00000000000000000001110101011101; // input=-3.373046875, output=0.229393208495
			11'd1888: out = 32'b00000000000000000001110111011001; // input=-3.376953125, output=0.233193533993
			11'd1889: out = 32'b00000000000000000001111001010110; // input=-3.380859375, output=0.236990301245
			11'd1890: out = 32'b00000000000000000001111011010010; // input=-3.384765625, output=0.240783452315
			11'd1891: out = 32'b00000000000000000001111101001110; // input=-3.388671875, output=0.244572929327
			11'd1892: out = 32'b00000000000000000001111111001010; // input=-3.392578125, output=0.248358674457
			11'd1893: out = 32'b00000000000000000010000001000110; // input=-3.396484375, output=0.252140629939
			11'd1894: out = 32'b00000000000000000010000011000010; // input=-3.400390625, output=0.255918738065
			11'd1895: out = 32'b00000000000000000010000100111110; // input=-3.404296875, output=0.259692941186
			11'd1896: out = 32'b00000000000000000010000110111001; // input=-3.408203125, output=0.263463181712
			11'd1897: out = 32'b00000000000000000010001000110101; // input=-3.412109375, output=0.267229402115
			11'd1898: out = 32'b00000000000000000010001010110000; // input=-3.416015625, output=0.270991544925
			11'd1899: out = 32'b00000000000000000010001100101011; // input=-3.419921875, output=0.274749552738
			11'd1900: out = 32'b00000000000000000010001110100110; // input=-3.423828125, output=0.27850336821
			11'd1901: out = 32'b00000000000000000010010000100001; // input=-3.427734375, output=0.282252934064
			11'd1902: out = 32'b00000000000000000010010010011100; // input=-3.431640625, output=0.285998193086
			11'd1903: out = 32'b00000000000000000010010100010110; // input=-3.435546875, output=0.289739088127
			11'd1904: out = 32'b00000000000000000010010110010001; // input=-3.439453125, output=0.293475562106
			11'd1905: out = 32'b00000000000000000010011000001011; // input=-3.443359375, output=0.297207558008
			11'd1906: out = 32'b00000000000000000010011010000101; // input=-3.447265625, output=0.30093501889
			11'd1907: out = 32'b00000000000000000010011011111111; // input=-3.451171875, output=0.304657887873
			11'd1908: out = 32'b00000000000000000010011101111001; // input=-3.455078125, output=0.308376108151
			11'd1909: out = 32'b00000000000000000010011111110011; // input=-3.458984375, output=0.31208962299
			11'd1910: out = 32'b00000000000000000010100001101100; // input=-3.462890625, output=0.315798375725
			11'd1911: out = 32'b00000000000000000010100011100101; // input=-3.466796875, output=0.319502309765
			11'd1912: out = 32'b00000000000000000010100101011111; // input=-3.470703125, output=0.323201368593
			11'd1913: out = 32'b00000000000000000010100111011000; // input=-3.474609375, output=0.326895495766
			11'd1914: out = 32'b00000000000000000010101001010001; // input=-3.478515625, output=0.330584634915
			11'd1915: out = 32'b00000000000000000010101011001001; // input=-3.482421875, output=0.33426872975
			11'd1916: out = 32'b00000000000000000010101101000010; // input=-3.486328125, output=0.337947724056
			11'd1917: out = 32'b00000000000000000010101110111010; // input=-3.490234375, output=0.341621561694
			11'd1918: out = 32'b00000000000000000010110000110010; // input=-3.494140625, output=0.345290186609
			11'd1919: out = 32'b00000000000000000010110010101011; // input=-3.498046875, output=0.348953542819
			11'd1920: out = 32'b00000000000000000010110100100010; // input=-3.501953125, output=0.352611574428
			11'd1921: out = 32'b00000000000000000010110110011010; // input=-3.505859375, output=0.356264225619
			11'd1922: out = 32'b00000000000000000010111000010010; // input=-3.509765625, output=0.359911440655
			11'd1923: out = 32'b00000000000000000010111010001001; // input=-3.513671875, output=0.363553163886
			11'd1924: out = 32'b00000000000000000010111100000000; // input=-3.517578125, output=0.367189339743
			11'd1925: out = 32'b00000000000000000010111101110111; // input=-3.521484375, output=0.370819912742
			11'd1926: out = 32'b00000000000000000010111111101110; // input=-3.525390625, output=0.374444827485
			11'd1927: out = 32'b00000000000000000011000001100100; // input=-3.529296875, output=0.378064028661
			11'd1928: out = 32'b00000000000000000011000011011011; // input=-3.533203125, output=0.381677461046
			11'd1929: out = 32'b00000000000000000011000101010001; // input=-3.537109375, output=0.385285069501
			11'd1930: out = 32'b00000000000000000011000111000111; // input=-3.541015625, output=0.388886798981
			11'd1931: out = 32'b00000000000000000011001000111101; // input=-3.544921875, output=0.392482594526
			11'd1932: out = 32'b00000000000000000011001010110011; // input=-3.548828125, output=0.39607240127
			11'd1933: out = 32'b00000000000000000011001100101000; // input=-3.552734375, output=0.399656164437
			11'd1934: out = 32'b00000000000000000011001110011101; // input=-3.556640625, output=0.403233829342
			11'd1935: out = 32'b00000000000000000011010000010010; // input=-3.560546875, output=0.406805341395
			11'd1936: out = 32'b00000000000000000011010010000111; // input=-3.564453125, output=0.410370646099
			11'd1937: out = 32'b00000000000000000011010011111100; // input=-3.568359375, output=0.413929689052
			11'd1938: out = 32'b00000000000000000011010101110000; // input=-3.572265625, output=0.417482415947
			11'd1939: out = 32'b00000000000000000011010111100100; // input=-3.576171875, output=0.421028772574
			11'd1940: out = 32'b00000000000000000011011001011000; // input=-3.580078125, output=0.42456870482
			11'd1941: out = 32'b00000000000000000011011011001100; // input=-3.583984375, output=0.42810215867
			11'd1942: out = 32'b00000000000000000011011101000000; // input=-3.587890625, output=0.431629080208
			11'd1943: out = 32'b00000000000000000011011110110011; // input=-3.591796875, output=0.435149415617
			11'd1944: out = 32'b00000000000000000011100000100110; // input=-3.595703125, output=0.438663111181
			11'd1945: out = 32'b00000000000000000011100010011001; // input=-3.599609375, output=0.442170113286
			11'd1946: out = 32'b00000000000000000011100100001100; // input=-3.603515625, output=0.445670368419
			11'd1947: out = 32'b00000000000000000011100101111110; // input=-3.607421875, output=0.44916382317
			11'd1948: out = 32'b00000000000000000011100111110000; // input=-3.611328125, output=0.452650424234
			11'd1949: out = 32'b00000000000000000011101001100010; // input=-3.615234375, output=0.45613011841
			11'd1950: out = 32'b00000000000000000011101011010100; // input=-3.619140625, output=0.459602852601
			11'd1951: out = 32'b00000000000000000011101101000110; // input=-3.623046875, output=0.463068573818
			11'd1952: out = 32'b00000000000000000011101110110111; // input=-3.626953125, output=0.466527229179
			11'd1953: out = 32'b00000000000000000011110000101000; // input=-3.630859375, output=0.469978765908
			11'd1954: out = 32'b00000000000000000011110010011001; // input=-3.634765625, output=0.473423131339
			11'd1955: out = 32'b00000000000000000011110100001010; // input=-3.638671875, output=0.476860272915
			11'd1956: out = 32'b00000000000000000011110101111010; // input=-3.642578125, output=0.480290138191
			11'd1957: out = 32'b00000000000000000011110111101010; // input=-3.646484375, output=0.48371267483
			11'd1958: out = 32'b00000000000000000011111001011010; // input=-3.650390625, output=0.487127830609
			11'd1959: out = 32'b00000000000000000011111011001010; // input=-3.654296875, output=0.490535553416
			11'd1960: out = 32'b00000000000000000011111100111001; // input=-3.658203125, output=0.493935791254
			11'd1961: out = 32'b00000000000000000011111110101000; // input=-3.662109375, output=0.49732849224
			11'd1962: out = 32'b00000000000000000100000000010111; // input=-3.666015625, output=0.500713604605
			11'd1963: out = 32'b00000000000000000100000010000110; // input=-3.669921875, output=0.504091076697
			11'd1964: out = 32'b00000000000000000100000011110100; // input=-3.673828125, output=0.507460856978
			11'd1965: out = 32'b00000000000000000100000101100011; // input=-3.677734375, output=0.510822894032
			11'd1966: out = 32'b00000000000000000100000111010001; // input=-3.681640625, output=0.514177136557
			11'd1967: out = 32'b00000000000000000100001000111110; // input=-3.685546875, output=0.517523533371
			11'd1968: out = 32'b00000000000000000100001010101100; // input=-3.689453125, output=0.520862033412
			11'd1969: out = 32'b00000000000000000100001100011001; // input=-3.693359375, output=0.52419258574
			11'd1970: out = 32'b00000000000000000100001110000110; // input=-3.697265625, output=0.527515139534
			11'd1971: out = 32'b00000000000000000100001111110010; // input=-3.701171875, output=0.530829644096
			11'd1972: out = 32'b00000000000000000100010001011111; // input=-3.705078125, output=0.534136048851
			11'd1973: out = 32'b00000000000000000100010011001011; // input=-3.708984375, output=0.537434303347
			11'd1974: out = 32'b00000000000000000100010100110110; // input=-3.712890625, output=0.540724357256
			11'd1975: out = 32'b00000000000000000100010110100010; // input=-3.716796875, output=0.544006160377
			11'd1976: out = 32'b00000000000000000100011000001101; // input=-3.720703125, output=0.547279662634
			11'd1977: out = 32'b00000000000000000100011001111000; // input=-3.724609375, output=0.550544814076
			11'd1978: out = 32'b00000000000000000100011011100011; // input=-3.728515625, output=0.553801564881
			11'd1979: out = 32'b00000000000000000100011101001101; // input=-3.732421875, output=0.557049865356
			11'd1980: out = 32'b00000000000000000100011110111000; // input=-3.736328125, output=0.560289665936
			11'd1981: out = 32'b00000000000000000100100000100001; // input=-3.740234375, output=0.563520917184
			11'd1982: out = 32'b00000000000000000100100010001011; // input=-3.744140625, output=0.566743569797
			11'd1983: out = 32'b00000000000000000100100011110100; // input=-3.748046875, output=0.5699575746
			11'd1984: out = 32'b00000000000000000100100101011101; // input=-3.751953125, output=0.573162882552
			11'd1985: out = 32'b00000000000000000100100111000110; // input=-3.755859375, output=0.576359444743
			11'd1986: out = 32'b00000000000000000100101000101111; // input=-3.759765625, output=0.579547212398
			11'd1987: out = 32'b00000000000000000100101010010111; // input=-3.763671875, output=0.582726136876
			11'd1988: out = 32'b00000000000000000100101011111111; // input=-3.767578125, output=0.58589616967
			11'd1989: out = 32'b00000000000000000100101101100110; // input=-3.771484375, output=0.58905726241
			11'd1990: out = 32'b00000000000000000100101111001110; // input=-3.775390625, output=0.59220936686
			11'd1991: out = 32'b00000000000000000100110000110101; // input=-3.779296875, output=0.595352434924
			11'd1992: out = 32'b00000000000000000100110010011011; // input=-3.783203125, output=0.598486418642
			11'd1993: out = 32'b00000000000000000100110100000010; // input=-3.787109375, output=0.601611270194
			11'd1994: out = 32'b00000000000000000100110101101000; // input=-3.791015625, output=0.604726941898
			11'd1995: out = 32'b00000000000000000100110111001101; // input=-3.794921875, output=0.607833386213
			11'd1996: out = 32'b00000000000000000100111000110011; // input=-3.798828125, output=0.610930555738
			11'd1997: out = 32'b00000000000000000100111010011000; // input=-3.802734375, output=0.614018403215
			11'd1998: out = 32'b00000000000000000100111011111101; // input=-3.806640625, output=0.617096881526
			11'd1999: out = 32'b00000000000000000100111101100010; // input=-3.810546875, output=0.620165943698
			11'd2000: out = 32'b00000000000000000100111111000110; // input=-3.814453125, output=0.623225542901
			11'd2001: out = 32'b00000000000000000101000000101010; // input=-3.818359375, output=0.626275632449
			11'd2002: out = 32'b00000000000000000101000010001101; // input=-3.822265625, output=0.629316165801
			11'd2003: out = 32'b00000000000000000101000011110001; // input=-3.826171875, output=0.632347096563
			11'd2004: out = 32'b00000000000000000101000101010100; // input=-3.830078125, output=0.635368378486
			11'd2005: out = 32'b00000000000000000101000110110110; // input=-3.833984375, output=0.638379965469
			11'd2006: out = 32'b00000000000000000101001000011001; // input=-3.837890625, output=0.64138181156
			11'd2007: out = 32'b00000000000000000101001001111011; // input=-3.841796875, output=0.644373870953
			11'd2008: out = 32'b00000000000000000101001011011101; // input=-3.845703125, output=0.647356097993
			11'd2009: out = 32'b00000000000000000101001100111110; // input=-3.849609375, output=0.650328447176
			11'd2010: out = 32'b00000000000000000101001110011111; // input=-3.853515625, output=0.653290873148
			11'd2011: out = 32'b00000000000000000101010000000000; // input=-3.857421875, output=0.656243330704
			11'd2012: out = 32'b00000000000000000101010001100000; // input=-3.861328125, output=0.659185774794
			11'd2013: out = 32'b00000000000000000101010011000000; // input=-3.865234375, output=0.662118160521
			11'd2014: out = 32'b00000000000000000101010100100000; // input=-3.869140625, output=0.665040443139
			11'd2015: out = 32'b00000000000000000101010101111111; // input=-3.873046875, output=0.667952578058
			11'd2016: out = 32'b00000000000000000101010111011111; // input=-3.876953125, output=0.670854520842
			11'd2017: out = 32'b00000000000000000101011000111101; // input=-3.880859375, output=0.673746227212
			11'd2018: out = 32'b00000000000000000101011010011100; // input=-3.884765625, output=0.676627653043
			11'd2019: out = 32'b00000000000000000101011011111010; // input=-3.888671875, output=0.679498754369
			11'd2020: out = 32'b00000000000000000101011101011000; // input=-3.892578125, output=0.68235948738
			11'd2021: out = 32'b00000000000000000101011110110101; // input=-3.896484375, output=0.685209808425
			11'd2022: out = 32'b00000000000000000101100000010010; // input=-3.900390625, output=0.688049674011
			11'd2023: out = 32'b00000000000000000101100001101111; // input=-3.904296875, output=0.690879040805
			11'd2024: out = 32'b00000000000000000101100011001011; // input=-3.908203125, output=0.693697865636
			11'd2025: out = 32'b00000000000000000101100100100111; // input=-3.912109375, output=0.69650610549
			11'd2026: out = 32'b00000000000000000101100110000011; // input=-3.916015625, output=0.699303717518
			11'd2027: out = 32'b00000000000000000101100111011110; // input=-3.919921875, output=0.702090659032
			11'd2028: out = 32'b00000000000000000101101000111001; // input=-3.923828125, output=0.704866887506
			11'd2029: out = 32'b00000000000000000101101010010100; // input=-3.927734375, output=0.707632360579
			11'd2030: out = 32'b00000000000000000101101011101110; // input=-3.931640625, output=0.710387036053
			11'd2031: out = 32'b00000000000000000101101101001000; // input=-3.935546875, output=0.713130871894
			11'd2032: out = 32'b00000000000000000101101110100001; // input=-3.939453125, output=0.715863826236
			11'd2033: out = 32'b00000000000000000101101111111011; // input=-3.943359375, output=0.718585857376
			11'd2034: out = 32'b00000000000000000101110001010011; // input=-3.947265625, output=0.72129692378
			11'd2035: out = 32'b00000000000000000101110010101100; // input=-3.951171875, output=0.723996984081
			11'd2036: out = 32'b00000000000000000101110100000100; // input=-3.955078125, output=0.726685997079
			11'd2037: out = 32'b00000000000000000101110101011100; // input=-3.958984375, output=0.729363921742
			11'd2038: out = 32'b00000000000000000101110110110011; // input=-3.962890625, output=0.732030717209
			11'd2039: out = 32'b00000000000000000101111000001010; // input=-3.966796875, output=0.734686342788
			11'd2040: out = 32'b00000000000000000101111001100001; // input=-3.970703125, output=0.737330757958
			11'd2041: out = 32'b00000000000000000101111010110111; // input=-3.974609375, output=0.739963922367
			11'd2042: out = 32'b00000000000000000101111100001101; // input=-3.978515625, output=0.742585795837
			11'd2043: out = 32'b00000000000000000101111101100011; // input=-3.982421875, output=0.745196338362
			11'd2044: out = 32'b00000000000000000101111110111000; // input=-3.986328125, output=0.747795510107
			11'd2045: out = 32'b00000000000000000110000000001101; // input=-3.990234375, output=0.750383271413
			11'd2046: out = 32'b00000000000000000110000001100001; // input=-3.994140625, output=0.752959582793
			11'd2047: out = 32'b00000000000000000110000010110101; // input=-3.998046875, output=0.755524404937
		endcase
	end
	converter U0 (a, index);

endmodule

module converter(a, index);
	input  [31:0] a;
	output [10:0] index;

	assign index[10]	= a[31];
	assign index[9:8]	= a[16:15];
	assign index[7:0]	= a[14:7];
endmodule
